----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:20:54 10/17/2016 
-- Design Name: 
-- Module Name:    Top - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
----------------------------------------------------------------------------------
-- VGA Colour Cycle
-- Michelle, 2015
----------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.ALL;
use IEEE.numeric_std.all;

entity VGATop is
  port(	clk50  : in std_logic;
		rst    : in std_logic;
		r      : out std_logic;
		g      : out std_logic;
		b      : out std_logic;
		hSync  : out std_logic;
		vSync  : out std_logic;
		UpButton : in std_logic;
		DownButton : in std_logic;
		rotary_a_in : in std_logic;
		rotary_b_in : in std_logic;
		--ROT_CENTER : in std_logic;
		fireButton : in std_logic);
		
end VGATop;


architecture RTL of VGATop is

-- Signals
signal clk25  : std_logic;
signal vidOn  : std_logic;
signal rgb    : std_logic_vector(2 downto 0);
signal row 	  : std_logic_vector(9 downto 0);
signal col    : std_logic_vector(9 downto 0);
signal rowInt : integer range 0 to 525;
signal colInt : integer range 0 to 800;
signal spaceShipX  : integer range 20 to 620;
signal clkCnt : std_logic_vector(24 downto 0);
signal clkTick : std_logic;
signal movementTick : std_logic;
signal scoreTick : std_logic;

signal score10000000000: integer range 0 to 10 := 0;
signal score1000000000: integer range 0 to 10 := 0;
signal score100000000: integer range 0 to 10 := 0;
signal score10000000: integer range 0 to 10 := 0;
signal score1000000: integer range 0 to 10 := 0;
signal score100000: integer range 0 to 10 := 0;
signal score10000: integer range 0 to 10 := 0;
signal score1000: integer range 0 to 10 := 0;
signal score100: integer range 0 to 10 := 0;
signal score10: integer range 0 to 10 := 0;

signal startdebounce : boolean := false;
signal debounceCounter : std_logic_vector(3 downto 0) := "1000";
signal fireSignal : std_logic;
signal bulletX : integer range 114 to 640; 
signal bulletY : integer range 0 to 480;

signal alien1_X : integer range 40 to 640; 
signal alien1_Y : integer range 50 to 420;
signal alien1_alive : std_logic;

signal alien2_X : integer range 40 to 640; 
signal alien2_Y : integer range 50 to 420;
signal alien2_alive : std_logic;

signal alien3_X : integer range 40 to 640; 
signal alien3_Y : integer range 50 to 420;
signal alien3_alive : std_logic;

signal alien4_X : integer range 40 to 640; 
signal alien4_Y : integer range 50 to 420;
signal alien4_alive : std_logic;

signal alien5_X : integer range 40 to 640; 
signal alien5_Y : integer range 50 to 420;
signal alien5_alive : std_logic;

signal rotary_in : std_logic_vector(1 downto 0) := "00";
signal rotary_q1 : std_logic;
signal rotary_q2 : std_logic;
signal rotary_left : std_logic;
signal rotary_event : std_logic;
signal delay_rotary_q1 : std_logic;

signal gameOver : std_logic;


type array_type_8x8 is array (7 downto 0) of unsigned (7 downto 0);


type array_type_16x16 is array (15 downto 0) of unsigned (15 downto 0);

Signal Score_0 : array_type_16x16;
Signal Score_1 : array_type_16x16;
Signal Score_2 : array_type_16x16;
Signal Score_3 : array_type_16x16;
Signal Score_4 : array_type_16x16;
Signal Score_5 : array_type_16x16;
Signal Score_6 : array_type_16x16;
Signal Score_7 : array_type_16x16;
Signal Score_8 : array_type_16x16;
Signal Score_9 : array_type_16x16;
Signal Score_Semi : array_type_16x16;
Signal Score_S : array_type_16x16;
Signal Score_C : array_type_16x16;
Signal Score_O : array_type_16x16;
Signal Score_R : array_type_16x16;
Signal Score_E : array_type_16x16;
Signal Score_Tracker10000000000 : array_type_16x16;
Signal Score_Tracker1000000000 : array_type_16x16;
Signal Score_Tracker100000000 : array_type_16x16;
Signal Score_Tracker10000000 : array_type_16x16;
Signal Score_Tracker1000000 : array_type_16x16;
Signal Score_Tracker100000 : array_type_16x16;
Signal Score_Tracker10000 : array_type_16x16;
Signal Score_Tracker1000 : array_type_16x16;
Signal Score_Tracker100 : array_type_16x16;
Signal Score_Tracker10 : array_type_16x16;
signal GameOver_V_W : array_type_16x16;
signal GameOver_A_W : array_type_16x16;
signal GameOver_G_W : array_type_16x16;
signal GameOver_M_W : array_type_16x16;

Signal Fire_Blast_1_R : array_type_16x16;
Signal Fire_Blast_1_G : array_type_16x16;
Signal Fire_Blast_1_B : array_type_16x16;

Signal Fire_Blast_2_R : array_type_16x16;
Signal Fire_Blast_2_G : array_type_16x16;
Signal Fire_Blast_2_B : array_type_16x16;


type array_type_32x32 is array (31 downto 0) of unsigned (31 downto 0);     -- only included once

signal Alien_1_R : array_type_32x32;
signal Alien_1_B : array_type_32x32;
signal Alien_1_G : array_type_32x32;

signal Alien_2_R : array_type_32x32;
signal Alien_2_G : array_type_32x32;
signal Alien_2_B : array_type_32x32;


type array_type_64x64 is array (63 downto 0) of unsigned (63 downto 0);

signal SpaceShip_Frame1_R : array_type_64x64;
signal SpaceShip_Frame1_G : array_type_64x64;
signal SpaceShip_Frame1_B : array_type_64x64;


signal SpaceShip_Frame2_R : array_type_64x64;
signal SpaceShip_Frame2_G : array_type_64x64;
signal SpaceShip_Frame2_B : array_type_64x64;

signal SpaceShip_Frame_Fire_R : array_type_64x64;
signal SpaceShip_Frame_Fire_G : array_type_64x64;
signal SpaceShip_Frame_Fire_B : array_type_64x64;


-- Components
component VGASync
	port(	clk	  :	in std_logic;
			rst	  :	in std_logic;
			hSync :	out std_logic;
			vSync :	out std_logic;
			row	  :	out std_logic_vector(9 downto 0);
			col	  :	out std_logic_vector(9 downto 0);
			vidOn :	out std_logic
	);
end component VGASync;
	
begin


Score_0(0) <= "0000011111100000";
Score_0(1) <= "0000011111100000";
Score_0(2) <= "0001100000011000";
Score_0(3) <= "0001100000011000";
Score_0(4) <= "0001100000011000";
Score_0(5) <= "0001100000011000";
Score_0(6) <= "0001100000011000";
Score_0(7) <= "0001100000011000";
Score_0(8) <= "0001100000011000";
Score_0(9) <= "0001100000011000";
Score_0(10) <= "0001100000011000";
Score_0(11) <= "0001100000011000";
Score_0(12) <= "0001100000011000";
Score_0(13) <= "0001100000011000";
Score_0(14) <= "0000011111100000";
Score_0(15) <= "0000011111100000";

Score_1(0) <= "0000000110000000";
Score_1(1) <= "0000001110000000";
Score_1(2) <= "0000011110000000";
Score_1(3) <= "0000000110000000";
Score_1(4) <= "0000000110000000";
Score_1(5) <= "0000000110000000";
Score_1(6) <= "0000000110000000";
Score_1(7) <= "0000000110000000";
Score_1(8) <= "0000000110000000";
Score_1(9) <= "0000000110000000";
Score_1(10) <= "0000000110000000";
Score_1(11) <= "0000000110000000";
Score_1(12) <= "0000000110000000";
Score_1(13) <= "0000000110000000";
Score_1(14) <= "0000011111100000";
Score_1(15) <= "0000011111100000";

Score_2(0) <= "0000111111110000";
Score_2(1) <= "0001111111111000";
Score_2(2) <= "0001100000011000";
Score_2(3) <= "0000000000011000";
Score_2(4) <= "0000000000011000";
Score_2(5) <= "0000000000011000";
Score_2(6) <= "0000000000110000";
Score_2(7) <= "0000000001100000";
Score_2(8) <= "0000000011000000";
Score_2(9) <= "0000000110000000";
Score_2(10) <= "0000001100000000";
Score_2(11) <= "0000011000000000";
Score_2(12) <= "0000110000000000";
Score_2(13) <= "0001111111111000";
Score_2(14) <= "0001111111111000";
Score_2(15) <= "0001111111111000";

Score_3(0) <= "0000011111100000";
Score_3(1) <= "0000111111110000";
Score_3(2) <= "0001100000111000";
Score_3(3) <= "0000000000011000";
Score_3(4) <= "0000000000011000";
Score_3(5) <= "0000000000011000";
Score_3(6) <= "0000000000111000";
Score_3(7) <= "0000000011110000";
Score_3(8) <= "0000000011110000";
Score_3(9) <= "0000000000111000";
Score_3(10) <= "0000000000011000";
Score_3(11) <= "0000000000011000";
Score_3(12) <= "0000000000011000";
Score_3(13) <= "0001100000111000";
Score_3(14) <= "0000111111110000";
Score_3(15) <= "0000011111100000";

Score_4(0) <= "0001100000011000";
Score_4(1) <= "0001100000011000";
Score_4(2) <= "0001100000011000";
Score_4(3) <= "0001100000011000";
Score_4(4) <= "0001100000011000";
Score_4(5) <= "0001100000011000";
Score_4(6) <= "0001100000011000";
Score_4(7) <= "0001111111111000";
Score_4(8) <= "0001111111111000";
Score_4(9) <= "0000000000011000";
Score_4(10) <= "0000000000011000";
Score_4(11) <= "0000000000011000";
Score_4(12) <= "0000000000011000";
Score_4(13) <= "0000000000011000";
Score_4(14) <= "0000000000011000";
Score_4(15) <= "0000000000011000";

Score_5(0) <= "0001111111111000";
Score_5(1) <= "0001111111111000";
Score_5(2) <= "0001100000000000";
Score_5(3) <= "0001100000000000";
Score_5(4) <= "0001100000000000";
Score_5(5) <= "0001100000000000";
Score_5(6) <= "0001100000000000";
Score_5(7) <= "0001111111100000";
Score_5(8) <= "0001111111110000";
Score_5(9) <= "0000000000111000";
Score_5(10) <= "0000000000011000";
Score_5(11) <= "0000000000011000";
Score_5(12) <= "0000000000011000";
Score_5(13) <= "0000000000111000";
Score_5(14) <= "0001111111110000";
Score_5(15) <= "0001111111100000";

Score_6(0) <= "0001111111111000";
Score_6(1) <= "0001111111111000";
Score_6(2) <= "0001100000000000";
Score_6(3) <= "0001100000000000";
Score_6(4) <= "0001100000000000";
Score_6(5) <= "0001100000000000";
Score_6(6) <= "0001100000000000";
Score_6(7) <= "0001100000000000";
Score_6(8) <= "0001111111111000";
Score_6(9) <= "0001111111111000";
Score_6(10) <= "0001110000111000";
Score_6(11) <= "0001110000111000";
Score_6(12) <= "0001110000111000";
Score_6(13) <= "0001110000111000";
Score_6(14) <= "0001111111111000";
Score_6(15) <= "0001111111111000";

Score_7(0) <= "0001111111111000";
Score_7(1) <= "0001111111111000";
Score_7(2) <= "0000000000011000";
Score_7(3) <= "0000000000011000";
Score_7(4) <= "0000000000110000";
Score_7(5) <= "0000000000110000";
Score_7(6) <= "0000000001100000";
Score_7(7) <= "0000000001100000";
Score_7(8) <= "0000000011000000";
Score_7(9) <= "0000000011000000";
Score_7(10) <= "0000000110000000";
Score_7(11) <= "0000000110000000";
Score_7(12) <= "0000001100000000";
Score_7(13) <= "0000001100000000";
Score_7(14) <= "0000011000000000";
Score_7(15) <= "0000011000000000";

Score_8(0) <= "0000011111100000";
Score_8(1) <= "0000011111100000";
Score_8(2) <= "0001100000011000";
Score_8(3) <= "0001100000011000";
Score_8(4) <= "0001100000011000";
Score_8(5) <= "0001100000011000";
Score_8(6) <= "0001100000011000";
Score_8(7) <= "0000011111100000";
Score_8(8) <= "0000011111100000";
Score_8(9) <= "0001100000011000";
Score_8(10) <= "0001100000011000";
Score_8(11) <= "0001100000011000";
Score_8(12) <= "0001100000011000";
Score_8(13) <= "0001100000011000";
Score_8(14) <= "0000011111100000";
Score_8(15) <= "0000011111100000";

Score_9(0) <= "0000111111110000";
Score_9(1) <= "0000110000110000";
Score_9(2) <= "0000110000110000";
Score_9(3) <= "0000110000110000";
Score_9(4) <= "0000110000110000";
Score_9(5) <= "0000110000110000";
Score_9(6) <= "0000111111110000";
Score_9(7) <= "0000111111110000";
Score_9(8) <= "0000000000110000";
Score_9(9) <= "0000000000110000";
Score_9(10) <= "0000000000110000";
Score_9(11) <= "0000000000110000";
Score_9(12) <= "0000000000110000";
Score_9(13) <= "0000000000110000";
Score_9(14) <= "0000111111110000";
Score_9(15) <= "0000111111110000";

Score_S(0) <= "0000011111111100";
Score_S(1) <= "0000111111111100";
Score_S(2) <= "0001110000000000";
Score_S(3) <= "0001100000000000";
Score_S(4) <= "0001100000000000";
Score_S(5) <= "0001100000000000";
Score_S(6) <= "0001110000000000";
Score_S(7) <= "0000111111110000";
Score_S(8) <= "0000011111111000";
Score_S(9) <= "0000000000001100";
Score_S(10) <= "0000000000001100";
Score_S(11) <= "0000000000001100";
Score_S(12) <= "0000000000001100";
Score_S(13) <= "0000000000011100";
Score_S(14) <= "0001111111111000";
Score_S(15) <= "0001111111110000";

Score_C(0) <= "0000111111111100";
Score_C(1) <= "0001111111111100";
Score_C(2) <= "0011100000000000";
Score_C(3) <= "0011000000000000";
Score_C(4) <= "0011000000000000";
Score_C(5) <= "0011000000000000";
Score_C(6) <= "0011000000000000";
Score_C(7) <= "0011000000000000";
Score_C(8) <= "0011000000000000";
Score_C(9) <= "0011000000000000";
Score_C(10) <= "0011000000000000";
Score_C(11) <= "0011000000000000";
Score_C(12) <= "0011000000000000";
Score_C(13) <= "0011100000000000";
Score_C(14) <= "0001111111111100";
Score_C(15) <= "0000111111111100";

Score_O(0) <= "0000111111110000";
Score_O(1) <= "0001111111111000";
Score_O(2) <= "0011100000011100";
Score_O(3) <= "0011000000001100";
Score_O(4) <= "0011000000001100";
Score_O(5) <= "0011000000001100";
Score_O(6) <= "0011000000001100";
Score_O(7) <= "0011000000001100";
Score_O(8) <= "0011000000001100";
Score_O(9) <= "0011000000001100";
Score_O(10) <= "0011000000001100";
Score_O(11) <= "0011000000001100";
Score_O(12) <= "0011000000001100";
Score_O(13) <= "0011100000011100";
Score_O(14) <= "0001111111111000";
Score_O(15) <= "0000111111110000";

Score_R(0) <= "0011111111110000";
Score_R(1) <= "0011111111111000";
Score_R(2) <= "0011000000011100";
Score_R(3) <= "0011000000001100";
Score_R(4) <= "0011000000001100";
Score_R(5) <= "0011000000011100";
Score_R(6) <= "0011000000111000";
Score_R(7) <= "0011111111110000";
Score_R(8) <= "0011111111110000";
Score_R(9) <= "0011000000111000";
Score_R(10) <= "0011000000011100";
Score_R(11) <= "0011000000001100";
Score_R(12) <= "0011000000001100";
Score_R(13) <= "0011000000001100";
Score_R(14) <= "0011000000001100";
Score_R(15) <= "0011000000001100";

Score_E(0) <= "0011111111111100";
Score_E(1) <= "0011111111111100";
Score_E(2) <= "0011000000000000";
Score_E(3) <= "0011000000000000";
Score_E(4) <= "0011000000000000";
Score_E(5) <= "0011000000000000";
Score_E(6) <= "0011000000000000";
Score_E(7) <= "0011111111110000";
Score_E(8) <= "0011111111110000";
Score_E(9) <= "0011000000000000";
Score_E(10) <= "0011000000000000";
Score_E(11) <= "0011000000000000";
Score_E(12) <= "0011000000000000";
Score_E(13) <= "0011000000000000";
Score_E(14) <= "0011111111111100";
Score_E(15) <= "0011111111111100";

Score_Semi(0) <= "0000000000000000";
Score_Semi(1) <= "0000000000000000";
Score_Semi(2) <= "0000001111000000";
Score_Semi(3) <= "0000001111000000";
Score_Semi(4) <= "0000001111000000";
Score_Semi(5) <= "0000001111000000";
Score_Semi(6) <= "0000000000000000";
Score_Semi(7) <= "0000000000000000";
Score_Semi(8) <= "0000000000000000";
Score_Semi(9) <= "0000000000000000";
Score_Semi(10) <= "0000001111000000";
Score_Semi(11) <= "0000001111000000";
Score_Semi(12) <= "0000001111000000";
Score_Semi(13) <= "0000001111000000";
Score_Semi(14) <= "0000000000000000";
Score_Semi(15) <= "0000000000000000";

GameOver_A_W(0) <= "0000000110000000";
GameOver_A_W(1) <= "0000001111000000";
GameOver_A_W(2) <= "0000011111100000";
GameOver_A_W(3) <= "0000111001110000";
GameOver_A_W(4) <= "0000110000110000";
GameOver_A_W(5) <= "0000110000110000";
GameOver_A_W(6) <= "0000110000110000";
GameOver_A_W(7) <= "0000110000110000";
GameOver_A_W(8) <= "0000110000110000";
GameOver_A_W(9) <= "0000111111110000";
GameOver_A_W(10) <= "0000111111110000";
GameOver_A_W(11) <= "0000110000110000";
GameOver_A_W(12) <= "0000110000110000";
GameOver_A_W(13) <= "0000110000110000";
GameOver_A_W(14) <= "0000110000110000";
GameOver_A_W(15) <= "0000110000110000";

GameOver_G_W(0) <= "0001111111100000";
GameOver_G_W(1) <= "0001111111100000";
GameOver_G_W(2) <= "0001100001100000";
GameOver_G_W(3) <= "0001100000000000";
GameOver_G_W(4) <= "0001100000000000";
GameOver_G_W(5) <= "0001100000000000";
GameOver_G_W(6) <= "0001100000000000";
GameOver_G_W(7) <= "0001100000000000";
GameOver_G_W(8) <= "0001100111111000";
GameOver_G_W(9) <= "0001100111111000";
GameOver_G_W(10) <= "0001100001100000";
GameOver_G_W(11) <= "0001100001100000";
GameOver_G_W(12) <= "0001100001100000";
GameOver_G_W(13) <= "0001100001100000";
GameOver_G_W(14) <= "0001111111100000";
GameOver_G_W(15) <= "0001111111100000";

GameOver_M_W(0) <= "0011000000001100";
GameOver_M_W(1) <= "0011100000011100";
GameOver_M_W(2) <= "0011110000111100";
GameOver_M_W(3) <= "0011111001111100";
GameOver_M_W(4) <= "0011011111101100";
GameOver_M_W(5) <= "0011001111001100";
GameOver_M_W(6) <= "0011000110001100";
GameOver_M_W(7) <= "0011000000001100";
GameOver_M_W(8) <= "0011000000001100";
GameOver_M_W(9) <= "0011000000001100";
GameOver_M_W(10) <= "0011000000001100";
GameOver_M_W(11) <= "0011000000001100";
GameOver_M_W(12) <= "0011000000001100";
GameOver_M_W(13) <= "0011000000001100";
GameOver_M_W(14) <= "0011000000001100";
GameOver_M_W(15) <= "0011000000001100";

GameOver_V_W(0) <= "0011000000001100";
GameOver_V_W(1) <= "0011000000001100";
GameOver_V_W(2) <= "0011100000011100";
GameOver_V_W(3) <= "0011100000011100";
GameOver_V_W(4) <= "0001110000111000";
GameOver_V_W(5) <= "0001110000111000";
GameOver_V_W(6) <= "0001110000111000";
GameOver_V_W(7) <= "0001110000111000";
GameOver_V_W(8) <= "0000111001110000";
GameOver_V_W(9) <= "0000111001110000";
GameOver_V_W(10) <= "0000111001110000";
GameOver_V_W(11) <= "0000011001100000";
GameOver_V_W(12) <= "0000011001100000";
GameOver_V_W(13) <= "0000011111100000";
GameOver_V_W(14) <= "0000001111000000";
GameOver_V_W(15) <= "0000000110000000";

Fire_Blast_1_R(0) <= "0000000000000000";
Fire_Blast_1_R(1) <= "0000000100100000";
Fire_Blast_1_R(2) <= "0000000010010000";
Fire_Blast_1_R(3) <= "0001000000001000";
Fire_Blast_1_R(4) <= "0100000111111100";
Fire_Blast_1_R(5) <= "0000001111001110";
Fire_Blast_1_R(6) <= "0000111100000011";
Fire_Blast_1_R(7) <= "0000011110000011";
Fire_Blast_1_R(8) <= "0100001111001110";
Fire_Blast_1_R(9) <= "0000100111111100";
Fire_Blast_1_R(10) <= "0000000000001000";
Fire_Blast_1_R(11) <= "0000000100010000";
Fire_Blast_1_R(12) <= "0000001000100000";
Fire_Blast_1_R(13) <= "0000000000000000";
Fire_Blast_1_R(14) <= "0000000000000000";
Fire_Blast_1_R(15) <= "0000000000000000";

Fire_Blast_1_G(0) <= "0000000000000000";
Fire_Blast_1_G(1) <= "0000000100100000";
Fire_Blast_1_G(2) <= "0000000010010000";
Fire_Blast_1_G(3) <= "0000000000001000";
Fire_Blast_1_G(4) <= "0000000000000100";
Fire_Blast_1_G(5) <= "0000000000000010";
Fire_Blast_1_G(6) <= "0000000000000001";
Fire_Blast_1_G(7) <= "0000000000000001";
Fire_Blast_1_G(8) <= "0000000000000010";
Fire_Blast_1_G(9) <= "0000000000000100";
Fire_Blast_1_G(10) <= "0000000000001000";
Fire_Blast_1_G(11) <= "0000000100010000";
Fire_Blast_1_G(12) <= "0000001000100000";
Fire_Blast_1_G(13) <= "0000000000000000";
Fire_Blast_1_G(14) <= "0000000000000000";
Fire_Blast_1_G(15) <= "0000000000000000";

Fire_Blast_1_B(0) <= "0000000000000000";
Fire_Blast_1_B(1) <= "0000000000000000";
Fire_Blast_1_B(2) <= "0000000000000000";
Fire_Blast_1_B(3) <= "0000000000000000";
Fire_Blast_1_B(4) <= "0000000000000000";
Fire_Blast_1_B(5) <= "0000000000110000";
Fire_Blast_1_B(6) <= "0000000011111100";
Fire_Blast_1_B(7) <= "0000000001111100";
Fire_Blast_1_B(8) <= "0000000000110000";
Fire_Blast_1_B(9) <= "0000000000000000";
Fire_Blast_1_B(10) <= "0000000000000000";
Fire_Blast_1_B(11) <= "0000000000000000";
Fire_Blast_1_B(12) <= "0000000000000000";
Fire_Blast_1_B(13) <= "0000000000000000";
Fire_Blast_1_B(14) <= "0000000000000000";
Fire_Blast_1_B(15) <= "0000000000000000";

Fire_Blast_2_R(0) <= "0000000000000000";
Fire_Blast_2_R(1) <= "0000000100100000";
Fire_Blast_2_R(2) <= "0000100010010000";
Fire_Blast_2_R(3) <= "0000010001001000";
Fire_Blast_2_R(4) <= "0001000111111100";
Fire_Blast_2_R(5) <= "1000001110001110";
Fire_Blast_2_R(6) <= "0010111000000011";
Fire_Blast_2_R(7) <= "0000011100000011";
Fire_Blast_2_R(8) <= "0001001111001110";
Fire_Blast_2_R(9) <= "1000000111111100";
Fire_Blast_2_R(10) <= "0000100001001000";
Fire_Blast_2_R(11) <= "0001000010010000";
Fire_Blast_2_R(12) <= "0000000100100000";
Fire_Blast_2_R(13) <= "0000000000000000";
Fire_Blast_2_R(14) <= "0000000000000000";
Fire_Blast_2_R(15) <= "0000000000000000";

Fire_Blast_2_G(0) <= "0000000000000000";
Fire_Blast_2_G(1) <= "0000000100100000";
Fire_Blast_2_G(2) <= "0000100010010000";
Fire_Blast_2_G(3) <= "0000010001001000";
Fire_Blast_2_G(4) <= "0000000000000100";
Fire_Blast_2_G(5) <= "0000000000000010";
Fire_Blast_2_G(6) <= "0000000000000001";
Fire_Blast_2_G(7) <= "0000000000000001";
Fire_Blast_2_G(8) <= "0000000000000010";
Fire_Blast_2_G(9) <= "0000000000000100";
Fire_Blast_2_G(10) <= "0000100001001000";
Fire_Blast_2_G(11) <= "0001000010010000";
Fire_Blast_2_G(12) <= "0000000100100000";
Fire_Blast_2_G(13) <= "0000000000000000";
Fire_Blast_2_G(14) <= "0000000000000000";
Fire_Blast_2_G(15) <= "0000000000000000";

Fire_Blast_2_B(0) <= "0000000000000000";
Fire_Blast_2_B(1) <= "0000000000000000";
Fire_Blast_2_B(2) <= "0000000000000000";
Fire_Blast_2_B(3) <= "0000000000000000";
Fire_Blast_2_B(4) <= "0000000000000000";
Fire_Blast_2_B(5) <= "0000000001110000";
Fire_Blast_2_B(6) <= "0000000111111100";
Fire_Blast_2_B(7) <= "0000000011111100";
Fire_Blast_2_B(8) <= "0000000000110000";
Fire_Blast_2_B(9) <= "0000000000000000";
Fire_Blast_2_B(10) <= "0000000000000000";
Fire_Blast_2_B(11) <= "0000000000000000";
Fire_Blast_2_B(12) <= "0000000000000000";
Fire_Blast_2_B(13) <= "0000000000000000";
Fire_Blast_2_B(14) <= "0000000000000000";
Fire_Blast_2_B(15) <= "0000000000000000";

Alien_1_R(0) <= "00000000000000000000000000000000";
Alien_1_R(1) <= "00000000000000000000000000000000";
Alien_1_R(2) <= "00000000000000000000000000000000";
Alien_1_R(3) <= "00000000000000000000000000000000";
Alien_1_R(4) <= "00000000000111111111100000000000";
Alien_1_R(5) <= "00000000001111111111110000000000";
Alien_1_R(6) <= "00000000010111111111101000000000";
Alien_1_R(7) <= "00000000101011111111010100000000";
Alien_1_R(8) <= "00000001110101111110101110000000";
Alien_1_R(9) <= "00000011111010111101011111000000";
Alien_1_R(10) <= "00000111111101100110111111100000";
Alien_1_R(11) <= "00001111111111100111111111110000";
Alien_1_R(12) <= "00000000000011100111000000000000";
Alien_1_R(13) <= "00000000000011000011000000000000";
Alien_1_R(14) <= "00001111111111011011111111110000";
Alien_1_R(15) <= "00001111111111011011111111110000";
Alien_1_R(16) <= "00001111111111011011111111110000";
Alien_1_R(17) <= "00000000000011000011000000000000";
Alien_1_R(18) <= "00000000000011100111000000000000";
Alien_1_R(19) <= "00001111111111100111111111110000";
Alien_1_R(20) <= "00001111111101100110111111110000";
Alien_1_R(21) <= "00000111111010111101011111100000";
Alien_1_R(22) <= "00000011110101111110101111000000";
Alien_1_R(23) <= "00000001101011111111010110000000";
Alien_1_R(24) <= "00000000010111111111101000000000";
Alien_1_R(25) <= "00000000001111111111110000000000";
Alien_1_R(26) <= "00000000001111111111110000000000";
Alien_1_R(27) <= "00000000000111111111100000000000";
Alien_1_R(28) <= "00000000000000000000000000000000";
Alien_1_R(29) <= "00000000000000000000000000000000";
Alien_1_R(30) <= "00000000000000000000000000000000";
Alien_1_R(31) <= "00000000000000000000000000000000";

Alien_1_G(0) <= "00000000000000000000000000000000";
Alien_1_G(1) <= "00000000000000000000000000000000";
Alien_1_G(2) <= "00000000000111111111100000000000";
Alien_1_G(3) <= "00000000001111111111110000000000";
Alien_1_G(4) <= "00000000011000011000011000000000";
Alien_1_G(5) <= "00000000110000011000001100000000";
Alien_1_G(6) <= "00000001101000011000010110000000";
Alien_1_G(7) <= "00000011000000011000000011000000";
Alien_1_G(8) <= "00000110001010011001010001100000";
Alien_1_G(9) <= "00001100000000111100000000110000";
Alien_1_G(10) <= "00011000000011111111000000011000";
Alien_1_G(11) <= "00110000000011111111000000001100";
Alien_1_G(12) <= "00111010101011111111010101011100";
Alien_1_G(13) <= "00110101010111111111101010101100";
Alien_1_G(14) <= "00110000000011100111000000001100";
Alien_1_G(15) <= "00110000000011100111000000001100";
Alien_1_G(16) <= "00110000000011100111000000001100";
Alien_1_G(17) <= "00110101010111111111101010101100";
Alien_1_G(18) <= "00111010101011111111010101011100";
Alien_1_G(19) <= "00110000000011111111000000001100";
Alien_1_G(20) <= "00110000000011111111000000001100";
Alien_1_G(21) <= "00011000000000111100000000011000";
Alien_1_G(22) <= "00001100001010011001010000110000";
Alien_1_G(23) <= "00000110000000011000000001100000";
Alien_1_G(24) <= "00000011101000011000010111000000";
Alien_1_G(25) <= "00000001100000011000000110000000";
Alien_1_G(26) <= "00000000110000011000001100000000";
Alien_1_G(27) <= "00000000011000011000011000000000";
Alien_1_G(28) <= "00000000001111111111110000000000";
Alien_1_G(29) <= "00000000000111111111100000000000";
Alien_1_G(30) <= "00000000000000000000000000000000";
Alien_1_G(31) <= "00000000000000000000000000000000";

Alien_1_B(0) <= "00000000001111111111110000000000";
Alien_1_B(1) <= "00000000001111111111110000000000";
Alien_1_B(2) <= "00000000011111111111111000000000";
Alien_1_B(3) <= "00000000111111111111111100000000";
Alien_1_B(4) <= "00000001111000000000011110000000";
Alien_1_B(5) <= "00000011110000000000001111000000";
Alien_1_B(6) <= "00000111100000000000000111100000";
Alien_1_B(7) <= "00001111010100000000101011110000";
Alien_1_B(8) <= "00011110000000000000000001111000";
Alien_1_B(9) <= "00111100000101000010100000111100";
Alien_1_B(10) <= "11111000000000000000000000011110";
Alien_1_B(11) <= "11110000000000100100000000001111";
Alien_1_B(12) <= "11110101010101100110101010101111";
Alien_1_B(13) <= "11111010101001000010010101011111";
Alien_1_B(14) <= "11110000000001000010000000001111";
Alien_1_B(15) <= "11110000000001000010000000001111";
Alien_1_B(16) <= "11110000000001000010000000001111";
Alien_1_B(17) <= "11111010101001000010010101011111";
Alien_1_B(18) <= "11110101010101100110101010101111";
Alien_1_B(19) <= "11110000000000100100000000001111";
Alien_1_B(20) <= "11110000000000000000000000001111";
Alien_1_B(21) <= "11111000000101000010100000011111";
Alien_1_B(22) <= "00111100000000000000000000111100";
Alien_1_B(23) <= "00011110010100000000101001111000";
Alien_1_B(24) <= "00001111000000000000000011110000";
Alien_1_B(25) <= "00000111110000000000001111100000";
Alien_1_B(26) <= "00000011110000000000001111000000";
Alien_1_B(27) <= "00000001111000000000011110000000";
Alien_1_B(28) <= "00000000111111111111111100000000";
Alien_1_B(29) <= "00000000011111111111111000000000";
Alien_1_B(30) <= "00000000001111111111110000000000";
Alien_1_B(31) <= "00000000001111111111110000000000";

Alien_2_R(0) <= "00000000000000000000000000000000";
Alien_2_R(1) <= "00000000000000000000000000000000";
Alien_2_R(2) <= "00000000000111111111100000000000";
Alien_2_R(3) <= "00000000001111111111110000000000";
Alien_2_R(4) <= "00000000011111100111111000000000";
Alien_2_R(5) <= "00000000111111100111111100000000";
Alien_2_R(6) <= "00000001110111100111101110000000";
Alien_2_R(7) <= "00000011101011100111010111000000";
Alien_2_R(8) <= "00000111110101100110101111100000";
Alien_2_R(9) <= "00001111111010000001011111110000";
Alien_2_R(10) <= "00011111111100000000111111111000";
Alien_2_R(11) <= "00111111111100100100111111111100";
Alien_2_R(12) <= "00110000000001100110000000001100";
Alien_2_R(13) <= "00110000000001000010000000001100";
Alien_2_R(14) <= "00111111111101011010111111111100";
Alien_2_R(15) <= "00111111111101011010111111111100";
Alien_2_R(16) <= "00111111111101011010111111111100";
Alien_2_R(17) <= "00110000000001000010000000001100";
Alien_2_R(18) <= "00110000000001100110000000001100";
Alien_2_R(19) <= "00111111111100100100111111111100";
Alien_2_R(20) <= "00111111111100000000111111111100";
Alien_2_R(21) <= "00011111111010000001011111111000";
Alien_2_R(22) <= "00001111110101100110101111110000";
Alien_2_R(23) <= "00000111101011100111010111100000";
Alien_2_R(24) <= "00000011010111100111101011000000";
Alien_2_R(25) <= "00000001101111100111110110000000";
Alien_2_R(26) <= "00000000111111100111111100000000";
Alien_2_R(27) <= "00000000011111100111111000000000";
Alien_2_R(28) <= "00000000001111111111110000000000";
Alien_2_R(29) <= "00000000000111111111100000000000";
Alien_2_R(30) <= "00000000000000000000000000000000";
Alien_2_R(31) <= "00000000000000000000000000000000";

Alien_2_G(0) <= "00000000000000000000000000000000";
Alien_2_G(1) <= "00000000000000000000000000000000";
Alien_2_G(2) <= "00000000000111111111100000000000";
Alien_2_G(3) <= "00000000001111111111110000000000";
Alien_2_G(4) <= "00000000011111111111111000000000";
Alien_2_G(5) <= "00000000111111111111111100000000";
Alien_2_G(6) <= "00000001110111111111101110000000";
Alien_2_G(7) <= "00000011111111111111111111000000";
Alien_2_G(8) <= "00000111110101111110101111100000";
Alien_2_G(9) <= "00001111111111111111111111110000";
Alien_2_G(10) <= "00011111111101111110111111111000";
Alien_2_G(11) <= "00111111111111011011111111111100";
Alien_2_G(12) <= "00110101010110011001101010101100";
Alien_2_G(13) <= "00111010101010111101010101011100";
Alien_2_G(14) <= "00111111111110111101111111111100";
Alien_2_G(15) <= "00111111111110111101111111111100";
Alien_2_G(16) <= "00111111111110111101111111111100";
Alien_2_G(17) <= "00111010101010111101010101011100";
Alien_2_G(18) <= "00110101010110011001101010101100";
Alien_2_G(19) <= "00111111111111011011111111111100";
Alien_2_G(20) <= "00111111111101111110111111111100";
Alien_2_G(21) <= "00011111111111111111111111111000";
Alien_2_G(22) <= "00001111110101111110101111110000";
Alien_2_G(23) <= "00000111111111111111111111100000";
Alien_2_G(24) <= "00000011010111111111101011000000";
Alien_2_G(25) <= "00000001111111111111111110000000";
Alien_2_G(26) <= "00000000111111111111111100000000";
Alien_2_G(27) <= "00000000011111111111111000000000";
Alien_2_G(28) <= "00000000001111111111110000000000";
Alien_2_G(29) <= "00000000000111111111100000000000";
Alien_2_G(30) <= "00000000000000000000000000000000";
Alien_2_G(31) <= "00000000000000000000000000000000";

Alien_2_B(0) <= "00000000001111111111110000000000";
Alien_2_B(1) <= "00000000001111111111110000000000";
Alien_2_B(2) <= "00000000011000000000011000000000";
Alien_2_B(3) <= "00000000110000000000001100000000";
Alien_2_B(4) <= "00000001100111111111100110000000";
Alien_2_B(5) <= "00000011001111111111110011000000";
Alien_2_B(6) <= "00000110011111111111111001100000";
Alien_2_B(7) <= "00001100101011111111010100110000";
Alien_2_B(8) <= "00011001111111111111111110011000";
Alien_2_B(9) <= "00110011111010111101011111001100";
Alien_2_B(10) <= "11100111111111100111111111100110";
Alien_2_B(11) <= "11001111111111000011111111110011";
Alien_2_B(12) <= "11001010101010000001010101010011";
Alien_2_B(13) <= "11000101010110000001101010100011";
Alien_2_B(14) <= "11001111111110011001111111110011";
Alien_2_B(15) <= "11001111111110011001111111110011";
Alien_2_B(16) <= "11001111111110011001111111110011";
Alien_2_B(17) <= "11000101010110000001101010100011";
Alien_2_B(18) <= "11001010101010000001010101010011";
Alien_2_B(19) <= "11001111111111000011111111110011";
Alien_2_B(20) <= "11001111111111100111111111110011";
Alien_2_B(21) <= "11100111111010111101011111100111";
Alien_2_B(22) <= "00110011111111111111111111001100";
Alien_2_B(23) <= "00011001101011111111010110011000";
Alien_2_B(24) <= "00001100111111111111111100110000";
Alien_2_B(25) <= "00000110001111111111110001100000";
Alien_2_B(26) <= "00000011001111111111110011000000";
Alien_2_B(27) <= "00000001100111111111100110000000";
Alien_2_B(28) <= "00000000110000000000001100000000";
Alien_2_B(29) <= "00000000011000000000011000000000";
Alien_2_B(30) <= "00000000001111111111110000000000";
Alien_2_B(31) <= "00000000001111111111110000000000";

SpaceShip_Frame1_R(0) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_R(1) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_R(2) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_R(3) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_R(4) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_R(5) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_R(6) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_R(7) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_R(8) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_R(9) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_R(10) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_R(11) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_R(12) <= "0000000000000000001111111100000000000000000000000000000000000000";
SpaceShip_Frame1_R(13) <= "0000000000000000001111111110000000000000000000000000000000000000";
SpaceShip_Frame1_R(14) <= "0000000000000000001111111111000000000000000000000000000000000000";
SpaceShip_Frame1_R(15) <= "0000000000000000001111111111100000000000000000000000000000000000";
SpaceShip_Frame1_R(16) <= "0000000000000000001111111111110000000000000000000000000000000000";
SpaceShip_Frame1_R(17) <= "0000000000000000001111111111111000000000000000000000000000000000";
SpaceShip_Frame1_R(18) <= "0000000000001111111111111111111100000000000000000000000000000000";
SpaceShip_Frame1_R(19) <= "0000000000001111111111111111111110000000000000000000000000000000";
SpaceShip_Frame1_R(20) <= "0000000000001111111111111111111111000000000000000000000000000000";
SpaceShip_Frame1_R(21) <= "0000000000001111111111111111111111100000000000000000000000000000";
SpaceShip_Frame1_R(22) <= "0000000000000111111111111111111111110000000000000000000000000000";
SpaceShip_Frame1_R(23) <= "0000000000000011111111111111111111111000000000000000000000000000";
SpaceShip_Frame1_R(24) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_R(25) <= "0000000000000000011111000000000000000000000000000000000000000000";
SpaceShip_Frame1_R(26) <= "0000000000000000000000000000000000010000000000000000000000000000";
SpaceShip_Frame1_R(27) <= "0000000000000000001110000000000000001000000000000000000000000000";
SpaceShip_Frame1_R(28) <= "0000000110000000000000000000000000000100000000000000000000000000";
SpaceShip_Frame1_R(29) <= "0000001111000000000100000000000000000010000000000000000000000000";
SpaceShip_Frame1_R(30) <= "0000011111100000000000000000000000000001000000000000000000000000";
SpaceShip_Frame1_R(31) <= "0001111111100000001110000000000000000000000000000000000000000000";
SpaceShip_Frame1_R(32) <= "0001111111100000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_R(33) <= "0000011111100000000100000000000000000001000000000000000000000000";
SpaceShip_Frame1_R(34) <= "0000001111000000000000000000000000000010000000000000000000000000";
SpaceShip_Frame1_R(35) <= "0000000110000000001110000000000000000100000000000000000000000000";
SpaceShip_Frame1_R(36) <= "0000000000000000000000000000000000001000000000000000000000000000";
SpaceShip_Frame1_R(37) <= "0000000000000000011111000000000000010000000000000000000000000000";
SpaceShip_Frame1_R(38) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_R(39) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_R(40) <= "0000000000000011111111111111111111111000000000000000000000000000";
SpaceShip_Frame1_R(41) <= "0000000000000111111111111111111111110000000000000000000000000000";
SpaceShip_Frame1_R(42) <= "0000000000001111111111111111111111100000000000000000000000000000";
SpaceShip_Frame1_R(43) <= "0000000000001111111111111111111111000000000000000000000000000000";
SpaceShip_Frame1_R(44) <= "0000000000001111111111111111111110000000000000000000000000000000";
SpaceShip_Frame1_R(45) <= "0000000000001111111111111111111100000000000000000000000000000000";
SpaceShip_Frame1_R(46) <= "0000000000000000001111111111111000000000000000000000000000000000";
SpaceShip_Frame1_R(47) <= "0000000000000000001111111111110000000000000000000000000000000000";
SpaceShip_Frame1_R(48) <= "0000000000000000001111111111100000000000000000000000000000000000";
SpaceShip_Frame1_R(49) <= "0000000000000000001111111111000000000000000000000000000000000000";
SpaceShip_Frame1_R(50) <= "0000000000000000001111111110000000000000000000000000000000000000";
SpaceShip_Frame1_R(51) <= "0000000000000000001111111100000000000000000000000000000000000000";
SpaceShip_Frame1_R(52) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_R(53) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_R(54) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_R(55) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_R(56) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_R(57) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_R(58) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_R(59) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_R(60) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_R(61) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_R(62) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_R(63) <= "0000000000000000000000000000000000000000000000000000000000000000";


SpaceShip_Frame1_G(0) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_G(1) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_G(2) <= "0000000000000001000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_G(3) <= "0000000000000001100000000000000000000000000000000000000000000000";
SpaceShip_Frame1_G(4) <= "0000000000000001110000000000000000000000000000000000000000000000";
SpaceShip_Frame1_G(5) <= "0000000000000001111000000000000000000000000000000000000000000000";
SpaceShip_Frame1_G(6) <= "0000000000000000111100000000000000000000000000000000000000000000";
SpaceShip_Frame1_G(7) <= "0000000000000000111110000000000000000000000000000000000000000000";
SpaceShip_Frame1_G(8) <= "0000000000000000011111000000000000000000000000000000000000000000";
SpaceShip_Frame1_G(9) <= "0000000000000000011111000000000000000000000000000000000000000000";
SpaceShip_Frame1_G(10) <= "0000000000000000011111110000000000000000000000000000000000000000";
SpaceShip_Frame1_G(11) <= "0000000000000000001111111000000000000000000000000000000000000000";
SpaceShip_Frame1_G(12) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_G(13) <= "0000000000000000001010101000000000000000000000000000000000000000";
SpaceShip_Frame1_G(14) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_G(15) <= "0000000000000000001111111111100011111110000000000000000000000000";
SpaceShip_Frame1_G(16) <= "0000000000000000000101010101010001111110000000000000000000000000";
SpaceShip_Frame1_G(17) <= "0000000000000000001111111111111000000000000000000000000000000000";
SpaceShip_Frame1_G(18) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_G(19) <= "0000000000001010101010101010101000000000000000000000000000000000";
SpaceShip_Frame1_G(20) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_G(21) <= "0000000000001111111111111111111111100000000000000000000000000000";
SpaceShip_Frame1_G(22) <= "0000000000000101010101010101010101110000000000000000000000000000";
SpaceShip_Frame1_G(23) <= "0000000000000011111111111111111111111000000000000000000000000000";
SpaceShip_Frame1_G(24) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_G(25) <= "0000000000000000000000000000111111111000000000000000000000000000";
SpaceShip_Frame1_G(26) <= "0000000000000000000000000001111111101100000000000000000000000000";
SpaceShip_Frame1_G(27) <= "0000000000000000000000000011111111110110000000000000000000000000";
SpaceShip_Frame1_G(28) <= "0000000000000000000000000111111111111011000000000000000000000000";
SpaceShip_Frame1_G(29) <= "0000000000000000000000001111111111111101100000000000000000000000";
SpaceShip_Frame1_G(30) <= "0000000000000000000000001111111111111110110000000000000000000000";
SpaceShip_Frame1_G(31) <= "0000000000000000000000001111111111111111111111111111111000000000";
SpaceShip_Frame1_G(32) <= "0000000000000000000000001111111111111111111111111111111000000000";
SpaceShip_Frame1_G(33) <= "0000000000000000000000001111111111111110110000000000000000000000";
SpaceShip_Frame1_G(34) <= "0000000000000000000000000111111111111101100000000000000000000000";
SpaceShip_Frame1_G(35) <= "0000000000000000000000000011111111111011000000000000000000000000";
SpaceShip_Frame1_G(36) <= "0000000000000000000000000001111111110110000000000000000000000000";
SpaceShip_Frame1_G(37) <= "0000000000000000000000000000111111101100000000000000000000000000";
SpaceShip_Frame1_G(38) <= "0000000000000000000000000000011111111000000000000000000000000000";
SpaceShip_Frame1_G(39) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_G(40) <= "0000000000000011111111111111111111111000000000000000000000000000";
SpaceShip_Frame1_G(41) <= "0000000000000101010101010101010101110000000000000000000000000000";
SpaceShip_Frame1_G(42) <= "0000000000001111111111111111111111100000000000000000000000000000";
SpaceShip_Frame1_G(43) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_G(44) <= "0000000000001010101010101010101000000000000000000000000000000000";
SpaceShip_Frame1_G(45) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_G(46) <= "0000000000000000001111111111111000000000000000000000000000000000";
SpaceShip_Frame1_G(47) <= "0000000000000000000101010101010001111110000000000000000000000000";
SpaceShip_Frame1_G(48) <= "0000000000000000001111111111100011111110000000000000000000000000";
SpaceShip_Frame1_G(49) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_G(50) <= "0000000000000000001010101000000000000000000000000000000000000000";
SpaceShip_Frame1_G(51) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_G(52) <= "0000000000000000001111111000000000000000000000000000000000000000";
SpaceShip_Frame1_G(53) <= "0000000000000000011111110000000000000000000000000000000000000000";
SpaceShip_Frame1_G(54) <= "0000000000000000011111100000000000000000000000000000000000000000";
SpaceShip_Frame1_G(55) <= "0000000000000000011111000000000000000000000000000000000000000000";
SpaceShip_Frame1_G(56) <= "0000000000000000111110000000000000000000000000000000000000000000";
SpaceShip_Frame1_G(57) <= "0000000000000000111100000000000000000000000000000000000000000000";
SpaceShip_Frame1_G(58) <= "0000000000000000111000000000000000000000000000000000000000000000";
SpaceShip_Frame1_G(59) <= "0000000000000001110000000000000000000000000000000000000000000000";
SpaceShip_Frame1_G(60) <= "0000000000000001100000000000000000000000000000000000000000000000";
SpaceShip_Frame1_G(61) <= "0000000000000001000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_G(62) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame1_G(63) <= "0000000000000000000000000000000000000000000000000000000000000000";

SpaceShip_Frame1_B(0) <= "0000000000001111100000000000000000000000000000000000000000000000";
SpaceShip_Frame1_B(1) <= "0000000000001111110000000000000000000000000000000000000000000000";
SpaceShip_Frame1_B(2) <= "0000000000001110111000000000000000000000000000000000000000000000";
SpaceShip_Frame1_B(3) <= "0000000000001110011100000000000000000000000000000000000000000000";
SpaceShip_Frame1_B(4) <= "0000000000000110001110000000000000000000000000000000000000000000";
SpaceShip_Frame1_B(5) <= "0000000000000110000111000000000000000000000000000000000000000000";
SpaceShip_Frame1_B(6) <= "0000000000000111000011100000000000000000000000000000000000000000";
SpaceShip_Frame1_B(7) <= "0000000000000011000001110000000000000000000000000000000000000000";
SpaceShip_Frame1_B(8) <= "0000000000000011100000111000000000000000000000000000000000000000";
SpaceShip_Frame1_B(9) <= "0000000000000011100000111100000000000000000000000000000000000000";
SpaceShip_Frame1_B(10) <= "0000000000000001100000001110000000000000000000000000000000000000";
SpaceShip_Frame1_B(11) <= "0000000000000001110000000111000000000000000000000000000000000000";
SpaceShip_Frame1_B(12) <= "0000011110000001110000000011100000000000000000000000000000000000";
SpaceShip_Frame1_B(13) <= "0000011111000000110000000001110000000000000000000000000000000000";
SpaceShip_Frame1_B(14) <= "0000011111100000110000000000111111111110000000000000000000000000";
SpaceShip_Frame1_B(15) <= "0000011111110000110000000000011100000001000000000000000000000000";
SpaceShip_Frame1_B(16) <= "0000011111111111110000000000001110000001000000000000000000000000";
SpaceShip_Frame1_B(17) <= "0000001111111111110000000000000111111110000000000000000000000000";
SpaceShip_Frame1_B(18) <= "0000000111110000000000000000000011100000000000000000000000000000";
SpaceShip_Frame1_B(19) <= "0000000011110000000000000000000001110000000000000000000000000000";
SpaceShip_Frame1_B(20) <= "0000000001110000000000000000000000111000000000000000000000000000";
SpaceShip_Frame1_B(21) <= "0000000000110000000000000000000000011100000000000000000000000000";
SpaceShip_Frame1_B(22) <= "0000000000011000000000000000000000001110000000000000000000000000";
SpaceShip_Frame1_B(23) <= "0000000000001100000000000000000000000111000000000000000000000000";
SpaceShip_Frame1_B(24) <= "0000000000000110000000000000000000000011100000000000000000000000";
SpaceShip_Frame1_B(25) <= "0000000000000110000000000000111111111001110000000000000000000000";
SpaceShip_Frame1_B(26) <= "0000000000000110000000000001111111111100111000000000000000000000";
SpaceShip_Frame1_B(27) <= "0000000000000110000000000011111111111110011100000100000000000000";
SpaceShip_Frame1_B(28) <= "0000000000000110000000000111111111111111001110000110000000000000";
SpaceShip_Frame1_B(29) <= "0000000000000110000000001111111111111111100111111111000000000000";
SpaceShip_Frame1_B(30) <= "0000000000001110000000001111111111111111110011111111111000000000";
SpaceShip_Frame1_B(31) <= "0000000000011110000000001111111111111111111111111111111100000000";
SpaceShip_Frame1_B(32) <= "0000000000011110000000001111111111111111111111111111111100000000";
SpaceShip_Frame1_B(33) <= "0000000000001110000000001111111111111111110011111111111000000000";
SpaceShip_Frame1_B(34) <= "0000000000000110000000000111111111111111100111111111000000000000";
SpaceShip_Frame1_B(35) <= "0000000000000110000000000011111111111111001110000110000000000000";
SpaceShip_Frame1_B(36) <= "0000000000000110000000000001111111111110011100000100000000000000";
SpaceShip_Frame1_B(37) <= "0000000000000110000000000000111111111100111000000000000000000000";
SpaceShip_Frame1_B(38) <= "0000000000000110000000000000011111111001110000000000000000000000";
SpaceShip_Frame1_B(39) <= "0000000000000110000000000000000000000011100000000000000000000000";
SpaceShip_Frame1_B(40) <= "0000000000001100000000000000000000000111000000000000000000000000";
SpaceShip_Frame1_B(41) <= "0000000000011000000000000000000000001110000000000000000000000000";
SpaceShip_Frame1_B(42) <= "0000000000110000000000000000000000011100000000000000000000000000";
SpaceShip_Frame1_B(43) <= "0000000001110000000000000000000000111000000000000000000000000000";
SpaceShip_Frame1_B(44) <= "0000000011110000000000000000000001110000000000000000000000000000";
SpaceShip_Frame1_B(45) <= "0000000111110000000000000000000011100000000000000000000000000000";
SpaceShip_Frame1_B(46) <= "0000001111111111110000000000000111111110000000000000000000000000";
SpaceShip_Frame1_B(47) <= "0000011111111111110000000000001110000001000000000000000000000000";
SpaceShip_Frame1_B(48) <= "0000011111110000110000000000011100000001000000000000000000000000";
SpaceShip_Frame1_B(49) <= "0000011111100000110000000000111111111110000000000000000000000000";
SpaceShip_Frame1_B(50) <= "0000011111000000110000000001110000000000000000000000000000000000";
SpaceShip_Frame1_B(51) <= "0000011110000001110000000011100000000000000000000000000000000000";
SpaceShip_Frame1_B(52) <= "0000000000000001110000000111000000000000000000000000000000000000";
SpaceShip_Frame1_B(53) <= "0000000000000001100000001110000000000000000000000000000000000000";
SpaceShip_Frame1_B(54) <= "0000000000000011100000011100000000000000000000000000000000000000";
SpaceShip_Frame1_B(55) <= "0000000000000011100000111000000000000000000000000000000000000000";
SpaceShip_Frame1_B(56) <= "0000000000000011000001110000000000000000000000000000000000000000";
SpaceShip_Frame1_B(57) <= "0000000000000111000011100000000000000000000000000000000000000000";
SpaceShip_Frame1_B(58) <= "0000000000000111000111000000000000000000000000000000000000000000";
SpaceShip_Frame1_B(59) <= "0000000000000110001110000000000000000000000000000000000000000000";
SpaceShip_Frame1_B(60) <= "0000000000001110011100000000000000000000000000000000000000000000";
SpaceShip_Frame1_B(61) <= "0000000000001110111000000000000000000000000000000000000000000000";
SpaceShip_Frame1_B(62) <= "0000000000001111110000000000000000000000000000000000000000000000";
SpaceShip_Frame1_B(63) <= "0000000000001111100000000000000000000000000000000000000000000000";


SpaceShip_Frame2_R(0) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_R(1) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_R(2) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_R(3) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_R(4) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_R(5) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_R(6) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_R(7) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_R(8) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_R(9) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_R(10) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_R(11) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_R(12) <= "0000000000000000001111111100000000000000000000000000000000000000";
SpaceShip_Frame2_R(13) <= "0000000000000000001111111110000000000000000000000000000000000000";
SpaceShip_Frame2_R(14) <= "0000000000000000001111111111000000000000000000000000000000000000";
SpaceShip_Frame2_R(15) <= "0000000000000000001111111111100000000000000000000000000000000000";
SpaceShip_Frame2_R(16) <= "0000000000000000001111111111110000000000000000000000000000000000";
SpaceShip_Frame2_R(17) <= "0000000000000000001111111111111000000000000000000000000000000000";
SpaceShip_Frame2_R(18) <= "0000000000001111111111111111111100000000000000000000000000000000";
SpaceShip_Frame2_R(19) <= "0000000000001111111111111111111110000000000000000000000000000000";
SpaceShip_Frame2_R(20) <= "0000000000001111111111111111111111000000000000000000000000000000";
SpaceShip_Frame2_R(21) <= "0000000000001111111111111111111111100000000000000000000000000000";
SpaceShip_Frame2_R(22) <= "0000000000000111111111111111111111110000000000000000000000000000";
SpaceShip_Frame2_R(23) <= "0000000000000011111111111111111111111000000000000000000000000000";
SpaceShip_Frame2_R(24) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_R(25) <= "0000000000000000011111000000000000000000000000000000000000000000";
SpaceShip_Frame2_R(26) <= "0000000000000000000000000000000000010000000000000000000000000000";
SpaceShip_Frame2_R(27) <= "0000000000000000001110000000000000001000000000000000000000000000";
SpaceShip_Frame2_R(28) <= "0000000000000000000000000000000000000100000000000000000000000000";
SpaceShip_Frame2_R(29) <= "0000000110000000000100000000000000000010000000000000000000000000";
SpaceShip_Frame2_R(30) <= "0100001111000000000000000000000000000001000000000000000000000000";
SpaceShip_Frame2_R(31) <= "0001011111100000001110000000000000000000000000000000000000000000";
SpaceShip_Frame2_R(32) <= "0000011111100000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_R(33) <= "0010001111000000000100000000000000000001000000000000000000000000";
SpaceShip_Frame2_R(34) <= "0000000110000000000000000000000000000010000000000000000000000000";
SpaceShip_Frame2_R(35) <= "0000000000000000001110000000000000000100000000000000000000000000";
SpaceShip_Frame2_R(36) <= "0000000000000000000000000000000000001000000000000000000000000000";
SpaceShip_Frame2_R(37) <= "0000000000000000011111000000000000010000000000000000000000000000";
SpaceShip_Frame2_R(38) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_R(39) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_R(40) <= "0000000000000011111111111111111111111000000000000000000000000000";
SpaceShip_Frame2_R(41) <= "0000000000000111111111111111111111110000000000000000000000000000";
SpaceShip_Frame2_R(42) <= "0000000000001111111111111111111111100000000000000000000000000000";
SpaceShip_Frame2_R(43) <= "0000000000001111111111111111111111000000000000000000000000000000";
SpaceShip_Frame2_R(44) <= "0000000000001111111111111111111110000000000000000000000000000000";
SpaceShip_Frame2_R(45) <= "0000000000001111111111111111111100000000000000000000000000000000";
SpaceShip_Frame2_R(46) <= "0000000000000000001111111111111000000000000000000000000000000000";
SpaceShip_Frame2_R(47) <= "0000000000000000001111111111110000000000000000000000000000000000";
SpaceShip_Frame2_R(48) <= "0000000000000000001111111111100000000000000000000000000000000000";
SpaceShip_Frame2_R(49) <= "0000000000000000001111111111000000000000000000000000000000000000";
SpaceShip_Frame2_R(50) <= "0000000000000000001111111110000000000000000000000000000000000000";
SpaceShip_Frame2_R(51) <= "0000000000000000001111111100000000000000000000000000000000000000";
SpaceShip_Frame2_R(52) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_R(53) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_R(54) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_R(55) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_R(56) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_R(57) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_R(58) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_R(59) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_R(60) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_R(61) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_R(62) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_R(63) <= "0000000000000000000000000000000000000000000000000000000000000000";


SpaceShip_Frame2_G(0) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_G(1) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_G(2) <= "0000000000000001000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_G(3) <= "0000000000000001100000000000000000000000000000000000000000000000";
SpaceShip_Frame2_G(4) <= "0000000000000001110000000000000000000000000000000000000000000000";
SpaceShip_Frame2_G(5) <= "0000000000000001111000000000000000000000000000000000000000000000";
SpaceShip_Frame2_G(6) <= "0000000000000000111100000000000000000000000000000000000000000000";
SpaceShip_Frame2_G(7) <= "0000000000000000111110000000000000000000000000000000000000000000";
SpaceShip_Frame2_G(8) <= "0000000000000000011111000000000000000000000000000000000000000000";
SpaceShip_Frame2_G(9) <= "0000000000000000011111000000000000000000000000000000000000000000";
SpaceShip_Frame2_G(10) <= "0000000000000000011111110000000000000000000000000000000000000000";
SpaceShip_Frame2_G(11) <= "0000000000000000001111111000000000000000000000000000000000000000";
SpaceShip_Frame2_G(12) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_G(13) <= "0000000000000000001010101000000000000000000000000000000000000000";
SpaceShip_Frame2_G(14) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_G(15) <= "0000000000000000001111111111100011111110000000000000000000000000";
SpaceShip_Frame2_G(16) <= "0000000000000000000101010101010001111110000000000000000000000000";
SpaceShip_Frame2_G(17) <= "0000000000000000001111111111111000000000000000000000000000000000";
SpaceShip_Frame2_G(18) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_G(19) <= "0000000000001010101010101010101000000000000000000000000000000000";
SpaceShip_Frame2_G(20) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_G(21) <= "0000000000001111111111111111111111100000000000000000000000000000";
SpaceShip_Frame2_G(22) <= "0000000000000101010101010101010101110000000000000000000000000000";
SpaceShip_Frame2_G(23) <= "0000000000000011111111111111111111111000000000000000000000000000";
SpaceShip_Frame2_G(24) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_G(25) <= "0000000000000000000000000000111111111000000000000000000000000000";
SpaceShip_Frame2_G(26) <= "0000000000000000000000000001111111101100000000000000000000000000";
SpaceShip_Frame2_G(27) <= "0000000000000000000000000011111111110110000000000000000000000000";
SpaceShip_Frame2_G(28) <= "0000000000000000000000000111111111111011000000000000000000000000";
SpaceShip_Frame2_G(29) <= "0000000000000000000000001111111111111101100000000000000000000000";
SpaceShip_Frame2_G(30) <= "0000000000000000000000001111111111111110110000000000000000000000";
SpaceShip_Frame2_G(31) <= "0000000000000000000000001111111111111111111111111111111000000000";
SpaceShip_Frame2_G(32) <= "0000000000000000000000001111111111111111111111111111111000000000";
SpaceShip_Frame2_G(33) <= "0000000000000000000000001111111111111110110000000000000000000000";
SpaceShip_Frame2_G(34) <= "0000000000000000000000000111111111111101100000000000000000000000";
SpaceShip_Frame2_G(35) <= "0000000000000000000000000011111111111011000000000000000000000000";
SpaceShip_Frame2_G(36) <= "0000000000000000000000000001111111110110000000000000000000000000";
SpaceShip_Frame2_G(37) <= "0000000000000000000000000000111111101100000000000000000000000000";
SpaceShip_Frame2_G(38) <= "0000000000000000000000000000011111111000000000000000000000000000";
SpaceShip_Frame2_G(39) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_G(40) <= "0000000000000011111111111111111111111000000000000000000000000000";
SpaceShip_Frame2_G(41) <= "0000000000000101010101010101010101110000000000000000000000000000";
SpaceShip_Frame2_G(42) <= "0000000000001111111111111111111111100000000000000000000000000000";
SpaceShip_Frame2_G(43) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_G(44) <= "0000000000001010101010101010101000000000000000000000000000000000";
SpaceShip_Frame2_G(45) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_G(46) <= "0000000000000000001111111111111000000000000000000000000000000000";
SpaceShip_Frame2_G(47) <= "0000000000000000000101010101010001111110000000000000000000000000";
SpaceShip_Frame2_G(48) <= "0000000000000000001111111111100011111110000000000000000000000000";
SpaceShip_Frame2_G(49) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_G(50) <= "0000000000000000001010101000000000000000000000000000000000000000";
SpaceShip_Frame2_G(51) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_G(52) <= "0000000000000000001111111000000000000000000000000000000000000000";
SpaceShip_Frame2_G(53) <= "0000000000000000011111110000000000000000000000000000000000000000";
SpaceShip_Frame2_G(54) <= "0000000000000000011111100000000000000000000000000000000000000000";
SpaceShip_Frame2_G(55) <= "0000000000000000011111000000000000000000000000000000000000000000";
SpaceShip_Frame2_G(56) <= "0000000000000000111110000000000000000000000000000000000000000000";
SpaceShip_Frame2_G(57) <= "0000000000000000111100000000000000000000000000000000000000000000";
SpaceShip_Frame2_G(58) <= "0000000000000000111000000000000000000000000000000000000000000000";
SpaceShip_Frame2_G(59) <= "0000000000000001110000000000000000000000000000000000000000000000";
SpaceShip_Frame2_G(60) <= "0000000000000001100000000000000000000000000000000000000000000000";
SpaceShip_Frame2_G(61) <= "0000000000000001000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_G(62) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame2_G(63) <= "0000000000000000000000000000000000000000000000000000000000000000";


SpaceShip_Frame2_B(0) <= "0000000000001111100000000000000000000000000000000000000000000000";
SpaceShip_Frame2_B(1) <= "0000000000001111110000000000000000000000000000000000000000000000";
SpaceShip_Frame2_B(2) <= "0000000000001110111000000000000000000000000000000000000000000000";
SpaceShip_Frame2_B(3) <= "0000000000001110011100000000000000000000000000000000000000000000";
SpaceShip_Frame2_B(4) <= "0000000000000110001110000000000000000000000000000000000000000000";
SpaceShip_Frame2_B(5) <= "0000000000000110000111000000000000000000000000000000000000000000";
SpaceShip_Frame2_B(6) <= "0000000000000111000011100000000000000000000000000000000000000000";
SpaceShip_Frame2_B(7) <= "0000000000000011000001110000000000000000000000000000000000000000";
SpaceShip_Frame2_B(8) <= "0000000000000011100000111000000000000000000000000000000000000000";
SpaceShip_Frame2_B(9) <= "0000000000000011100000111100000000000000000000000000000000000000";
SpaceShip_Frame2_B(10) <= "0000000000000001100000001110000000000000000000000000000000000000";
SpaceShip_Frame2_B(11) <= "0000000000000001110000000111000000000000000000000000000000000000";
SpaceShip_Frame2_B(12) <= "0000011110000001110000000011100000000000000000000000000000000000";
SpaceShip_Frame2_B(13) <= "0000011111000000110000000001110000000000000000000000000000000000";
SpaceShip_Frame2_B(14) <= "0000011111100000110000000000111111111110000000000000000000000000";
SpaceShip_Frame2_B(15) <= "0000011111110000110000000000011100000001000000000000000000000000";
SpaceShip_Frame2_B(16) <= "0000011111111111110000000000001110000001000000000000000000000000";
SpaceShip_Frame2_B(17) <= "0000001111111111110000000000000111111110000000000000000000000000";
SpaceShip_Frame2_B(18) <= "0000000111110000000000000000000011100000000000000000000000000000";
SpaceShip_Frame2_B(19) <= "0000000011110000000000000000000001110000000000000000000000000000";
SpaceShip_Frame2_B(20) <= "0000000001110000000000000000000000111000000000000000000000000000";
SpaceShip_Frame2_B(21) <= "0000000000110000000000000000000000011100000000000000000000000000";
SpaceShip_Frame2_B(22) <= "0000000000011000000000000000000000001110000000000000000000000000";
SpaceShip_Frame2_B(23) <= "0000000000001100000000000000000000000111000000000000000000000000";
SpaceShip_Frame2_B(24) <= "0000000000000110000000000000000000000011100000000000000000000000";
SpaceShip_Frame2_B(25) <= "0000000000000110000000000000111111111001110000000000000000000000";
SpaceShip_Frame2_B(26) <= "0000000000000110000000000001111111111100111000000000000000000000";
SpaceShip_Frame2_B(27) <= "0000000000000110000000000011111111111110011100000100000000000000";
SpaceShip_Frame2_B(28) <= "0000000000000110000000000111111111111111001110000110000000000000";
SpaceShip_Frame2_B(29) <= "0000000000000110000000001111111111111111100111111111000000000000";
SpaceShip_Frame2_B(30) <= "0000000000001110000000001111111111111111110011111111111000000000";
SpaceShip_Frame2_B(31) <= "0000000000011110000000001111111111111111111111111111111100000000";
SpaceShip_Frame2_B(32) <= "0000000000011110000000001111111111111111111111111111111100000000";
SpaceShip_Frame2_B(33) <= "0000000000001110000000001111111111111111110011111111111000000000";
SpaceShip_Frame2_B(34) <= "0000000000000110000000000111111111111111100111111111000000000000";
SpaceShip_Frame2_B(35) <= "0000000000000110000000000011111111111111001110000110000000000000";
SpaceShip_Frame2_B(36) <= "0000000000000110000000000001111111111110011100000100000000000000";
SpaceShip_Frame2_B(37) <= "0000000000000110000000000000111111111100111000000000000000000000";
SpaceShip_Frame2_B(38) <= "0000000000000110000000000000011111111001110000000000000000000000";
SpaceShip_Frame2_B(39) <= "0000000000000110000000000000000000000011100000000000000000000000";
SpaceShip_Frame2_B(40) <= "0000000000001100000000000000000000000111000000000000000000000000";
SpaceShip_Frame2_B(41) <= "0000000000011000000000000000000000001110000000000000000000000000";
SpaceShip_Frame2_B(42) <= "0000000000110000000000000000000000011100000000000000000000000000";
SpaceShip_Frame2_B(43) <= "0000000001110000000000000000000000111000000000000000000000000000";
SpaceShip_Frame2_B(44) <= "0000000011110000000000000000000001110000000000000000000000000000";
SpaceShip_Frame2_B(45) <= "0000000111110000000000000000000011100000000000000000000000000000";
SpaceShip_Frame2_B(46) <= "0000001111111111110000000000000111111110000000000000000000000000";
SpaceShip_Frame2_B(47) <= "0000011111111111110000000000001110000001000000000000000000000000";
SpaceShip_Frame2_B(48) <= "0000011111110000110000000000011100000001000000000000000000000000";
SpaceShip_Frame2_B(49) <= "0000011111100000110000000000111111111110000000000000000000000000";
SpaceShip_Frame2_B(50) <= "0000011111000000110000000001110000000000000000000000000000000000";
SpaceShip_Frame2_B(51) <= "0000011110000001110000000011100000000000000000000000000000000000";
SpaceShip_Frame2_B(52) <= "0000000000000001110000000111000000000000000000000000000000000000";
SpaceShip_Frame2_B(53) <= "0000000000000001100000001110000000000000000000000000000000000000";
SpaceShip_Frame2_B(54) <= "0000000000000011100000011100000000000000000000000000000000000000";
SpaceShip_Frame2_B(55) <= "0000000000000011100000111000000000000000000000000000000000000000";
SpaceShip_Frame2_B(56) <= "0000000000000011000001110000000000000000000000000000000000000000";
SpaceShip_Frame2_B(57) <= "0000000000000111000011100000000000000000000000000000000000000000";
SpaceShip_Frame2_B(58) <= "0000000000000111000111000000000000000000000000000000000000000000";
SpaceShip_Frame2_B(59) <= "0000000000000110001110000000000000000000000000000000000000000000";
SpaceShip_Frame2_B(60) <= "0000000000001110011100000000000000000000000000000000000000000000";
SpaceShip_Frame2_B(61) <= "0000000000001110111000000000000000000000000000000000000000000000";
SpaceShip_Frame2_B(62) <= "0000000000001111110000000000000000000000000000000000000000000000";
SpaceShip_Frame2_B(63) <= "0000000000001111100000000000000000000000000000000000000000000000";

SpaceShip_Frame_Fire_R(0) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(1) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(2) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(3) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(4) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(5) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(6) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(7) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(8) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(9) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(10) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(11) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(12) <= "0000000000000000001111111100000000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(13) <= "0000000000000000001111111110000000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(14) <= "0000000000000000001111111111000000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(15) <= "0000000000000000001111111111100000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(16) <= "0000000000000000001111111111110000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(17) <= "0000000000000000001111111111111000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(18) <= "0000000000001111111111111111111100000000000000000000000000000000";
SpaceShip_Frame_Fire_R(19) <= "0000000000001111111111111111111110000000000000000000000000000000";
SpaceShip_Frame_Fire_R(20) <= "0000000000001111111111111111111111000000000000000000000000000000";
SpaceShip_Frame_Fire_R(21) <= "0000000000001111111111111111111111100000000000000000000000000000";
SpaceShip_Frame_Fire_R(22) <= "0000000000000111111111111111111111110000000000000000000000000000";
SpaceShip_Frame_Fire_R(23) <= "0000000000000011111111111111111111111000000000000000000000000000";
SpaceShip_Frame_Fire_R(24) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(25) <= "0000000000000000011111000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(26) <= "0000000000000000000000000000000000010000000000000000000000011000";
SpaceShip_Frame_Fire_R(27) <= "0000000000000000001110000000000000001000000000000000000001100000";
SpaceShip_Frame_Fire_R(28) <= "0000000000000000000000000000000000000100000000000000000000000000";
SpaceShip_Frame_Fire_R(29) <= "0000000110000000000100000000000000000010000000000000000110110000";
SpaceShip_Frame_Fire_R(30) <= "0100001111000000000000000000000000000001000000000000000000000000";
SpaceShip_Frame_Fire_R(31) <= "0001011111100000001110000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(32) <= "0000011111100000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(33) <= "0010001111000000000100000000000000000001000000000000000000000000";
SpaceShip_Frame_Fire_R(34) <= "0000000110000000000000000000000000000010000000000000000110110000";
SpaceShip_Frame_Fire_R(35) <= "0000000000000000001110000000000000000100000000000000000000000000";
SpaceShip_Frame_Fire_R(36) <= "0000000000000000000000000000000000001000000000000000000001100000";
SpaceShip_Frame_Fire_R(37) <= "0000000000000000011111000000000000010000000000000000000000011000";
SpaceShip_Frame_Fire_R(38) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(39) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(40) <= "0000000000000011111111111111111111111000000000000000000000000000";
SpaceShip_Frame_Fire_R(41) <= "0000000000000111111111111111111111110000000000000000000000000000";
SpaceShip_Frame_Fire_R(42) <= "0000000000001111111111111111111111100000000000000000000000000000";
SpaceShip_Frame_Fire_R(43) <= "0000000000001111111111111111111111000000000000000000000000000000";
SpaceShip_Frame_Fire_R(44) <= "0000000000001111111111111111111110000000000000000000000000000000";
SpaceShip_Frame_Fire_R(45) <= "0000000000001111111111111111111100000000000000000000000000000000";
SpaceShip_Frame_Fire_R(46) <= "0000000000000000001111111111111000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(47) <= "0000000000000000001111111111110000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(48) <= "0000000000000000001111111111100000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(49) <= "0000000000000000001111111111000000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(50) <= "0000000000000000001111111110000000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(51) <= "0000000000000000001111111100000000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(52) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(53) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(54) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(55) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(56) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(57) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(58) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(59) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(60) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(61) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(62) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_R(63) <= "0000000000000000000000000000000000000000000000000000000000000000";


SpaceShip_Frame_Fire_G(0) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(1) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(2) <= "0000000000000001000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(3) <= "0000000000000001100000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(4) <= "0000000000000001110000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(5) <= "0000000000000001111000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(6) <= "0000000000000000111100000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(7) <= "0000000000000000111110000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(8) <= "0000000000000000011111000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(9) <= "0000000000000000011111100000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(10) <= "0000000000000000011111110000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(11) <= "0000000000000000001111111000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(12) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(13) <= "0000000000000000001010101000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(14) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(15) <= "0000000000000000001111111111100011111110000000000000000000000000";
SpaceShip_Frame_Fire_G(16) <= "0000000000000000000101010101010001111110000000000000000000000000";
SpaceShip_Frame_Fire_G(17) <= "0000000000000000001111111111111000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(18) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(19) <= "0000000000001010101010101010101000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(20) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(21) <= "0000000000001111111111111111111111100000000000000000000000000000";
SpaceShip_Frame_Fire_G(22) <= "0000000000000101010101010101010101110000000000000000000000000000";
SpaceShip_Frame_Fire_G(23) <= "0000000000000011111111111111111111111000000000000000000000000000";
SpaceShip_Frame_Fire_G(24) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(25) <= "0000000000000000000000000000111111111000000000000000000000000000";
SpaceShip_Frame_Fire_G(26) <= "0000000000000000000000000001111111101100000000000000000000010000";
SpaceShip_Frame_Fire_G(27) <= "0000000000000000000000000011111111110110000000000000000001000000";
SpaceShip_Frame_Fire_G(28) <= "0000000000000000000000000111111111111011000000000000000000000000";
SpaceShip_Frame_Fire_G(29) <= "0000000000000000000000001111111111111101100000000000000100100000";
SpaceShip_Frame_Fire_G(30) <= "0000000000000000000000001111111111111110110000000000000000000000";
SpaceShip_Frame_Fire_G(31) <= "0000000000000000000000001111111111111111111111111111111000000000";
SpaceShip_Frame_Fire_G(32) <= "0000000000000000000000001111111111111111111111111111111000000000";
SpaceShip_Frame_Fire_G(33) <= "0000000000000000000000001111111111111110110000000000000000000000";
SpaceShip_Frame_Fire_G(34) <= "0000000000000000000000000111111111111101100000000000000100100000";
SpaceShip_Frame_Fire_G(35) <= "0000000000000000000000000011111111111011000000000000000000000000";
SpaceShip_Frame_Fire_G(36) <= "0000000000000000000000000001111111110110000000000000000001000000";
SpaceShip_Frame_Fire_G(37) <= "0000000000000000000000000000111111101100000000000000000000010000";
SpaceShip_Frame_Fire_G(38) <= "0000000000000000000000000000011111111000000000000000000000000000";
SpaceShip_Frame_Fire_G(39) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(40) <= "0000000000000011111111111111111111111000000000000000000000000000";
SpaceShip_Frame_Fire_G(41) <= "0000000000000101010101010101010101110000000000000000000000000000";
SpaceShip_Frame_Fire_G(42) <= "0000000000001111111111111111111111100000000000000000000000000000";
SpaceShip_Frame_Fire_G(43) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(44) <= "0000000000001010101010101010101000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(45) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(46) <= "0000000000000000001111111111111000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(47) <= "0000000000000000000101010101010001111110000000000000000000000000";
SpaceShip_Frame_Fire_G(48) <= "0000000000000000001111111111100011111110000000000000000000000000";
SpaceShip_Frame_Fire_G(49) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(50) <= "0000000000000000001010101000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(51) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(52) <= "0000000000000000001111111000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(53) <= "0000000000000000011111110000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(54) <= "0000000000000000011111100000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(55) <= "0000000000000000011111000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(56) <= "0000000000000000111110000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(57) <= "0000000000000000111100000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(58) <= "0000000000000000111000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(59) <= "0000000000000001110000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(60) <= "0000000000000001100000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(61) <= "0000000000000001000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(62) <= "0000000000000000000000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_G(63) <= "0000000000000000000000000000000000000000000000000000000000000000";


SpaceShip_Frame_Fire_B(0) <= "0000000000001111100000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_B(1) <= "0000000000001111110000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_B(2) <= "0000000000001110111000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_B(3) <= "0000000000001110011100000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_B(4) <= "0000000000000110001110000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_B(5) <= "0000000000000110000111000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_B(6) <= "0000000000000111000011100000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_B(7) <= "0000000000000011000001110000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_B(8) <= "0000000000000011100000111000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_B(9) <= "0000000000000011100000011100000000000000000000000000000000000000";
SpaceShip_Frame_Fire_B(10) <= "0000000000000001100000001110000000000000000000000000000000000000";
SpaceShip_Frame_Fire_B(11) <= "0000000000000001110000000111000000000000000000000000000000000000";
SpaceShip_Frame_Fire_B(12) <= "0000011110000001110000000011100000000000000000000000000000000000";
SpaceShip_Frame_Fire_B(13) <= "0000011111000000110000000001110000000000000000000000000000000000";
SpaceShip_Frame_Fire_B(14) <= "0000011111100000110000000000111111111110000000000000000000000000";
SpaceShip_Frame_Fire_B(15) <= "0000011111110000110000000000011100000001000000000000000000000000";
SpaceShip_Frame_Fire_B(16) <= "0000011111111111110000000000001110000001000000000000000000000000";
SpaceShip_Frame_Fire_B(17) <= "0000001111111111110000000000000111111110000000000000000000000000";
SpaceShip_Frame_Fire_B(18) <= "0000000111110000000000000000000011100000000000000000000000000000";
SpaceShip_Frame_Fire_B(19) <= "0000000011110000000000000000000001110000000000000000000000000000";
SpaceShip_Frame_Fire_B(20) <= "0000000001110000000000000000000000111000000000000000000000000000";
SpaceShip_Frame_Fire_B(21) <= "0000000000110000000000000000000000011100000000000000000000000000";
SpaceShip_Frame_Fire_B(22) <= "0000000000011000000000000000000000001110000000000000000000000000";
SpaceShip_Frame_Fire_B(23) <= "0000000000001100000000000000000000000111000000000000000000000000";
SpaceShip_Frame_Fire_B(24) <= "0000000000000110000000000000000000000011100000000000000000000000";
SpaceShip_Frame_Fire_B(25) <= "0000000000000110000000000000111111111001110000000000000000000000";
SpaceShip_Frame_Fire_B(26) <= "0000000000000110000000000001111111111100111000000000000000000000";
SpaceShip_Frame_Fire_B(27) <= "0000000000000110000000000011111111111110011100000100000000000000";
SpaceShip_Frame_Fire_B(28) <= "0000000000000110000000000111111111111111001110000110000000000000";
SpaceShip_Frame_Fire_B(29) <= "0000000000000110000000001111111111111111100111111111000000000000";
SpaceShip_Frame_Fire_B(30) <= "0000000000001110000000001111111111111111110011111111111000000000";
SpaceShip_Frame_Fire_B(31) <= "0000000000011110000000001111111111111111111111111111111100000000";
SpaceShip_Frame_Fire_B(32) <= "0000000000011110000000001111111111111111111111111111111100000000";
SpaceShip_Frame_Fire_B(33) <= "0000000000001110000000001111111111111111110011111111111000000000";
SpaceShip_Frame_Fire_B(34) <= "0000000000000110000000000111111111111111100111111111000000000000";
SpaceShip_Frame_Fire_B(35) <= "0000000000000110000000000011111111111111001110000110000000000000";
SpaceShip_Frame_Fire_B(36) <= "0000000000000110000000000001111111111110011100000100000000000000";
SpaceShip_Frame_Fire_B(37) <= "0000000000000110000000000000111111111100111000000000000000000000";
SpaceShip_Frame_Fire_B(38) <= "0000000000000110000000000000011111111001110000000000000000000000";
SpaceShip_Frame_Fire_B(39) <= "0000000000000110000000000000000000000011100000000000000000000000";
SpaceShip_Frame_Fire_B(40) <= "0000000000001100000000000000000000000111000000000000000000000000";
SpaceShip_Frame_Fire_B(41) <= "0000000000011000000000000000000000001110000000000000000000000000";
SpaceShip_Frame_Fire_B(42) <= "0000000000110000000000000000000000011100000000000000000000000000";
SpaceShip_Frame_Fire_B(43) <= "0000000001110000000000000000000000111000000000000000000000000000";
SpaceShip_Frame_Fire_B(44) <= "0000000011110000000000000000000001110000000000000000000000000000";
SpaceShip_Frame_Fire_B(45) <= "0000000111110000000000000000000011100000000000000000000000000000";
SpaceShip_Frame_Fire_B(46) <= "0000001111111111110000000000000111111110000000000000000000000000";
SpaceShip_Frame_Fire_B(47) <= "0000011111111111110000000000001110000001000000000000000000000000";
SpaceShip_Frame_Fire_B(48) <= "0000011111110000110000000000011100000001000000000000000000000000";
SpaceShip_Frame_Fire_B(49) <= "0000011111100000110000000000111111111110000000000000000000000000";
SpaceShip_Frame_Fire_B(50) <= "0000011111000000110000000001110000000000000000000000000000000000";
SpaceShip_Frame_Fire_B(51) <= "0000011110000001110000000011100000000000000000000000000000000000";
SpaceShip_Frame_Fire_B(52) <= "0000000000000001110000000111000000000000000000000000000000000000";
SpaceShip_Frame_Fire_B(53) <= "0000000000000001100000001110000000000000000000000000000000000000";
SpaceShip_Frame_Fire_B(54) <= "0000000000000011100000011100000000000000000000000000000000000000";
SpaceShip_Frame_Fire_B(55) <= "0000000000000011100000111000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_B(56) <= "0000000000000011000001110000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_B(57) <= "0000000000000111000011100000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_B(58) <= "0000000000000111000111000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_B(59) <= "0000000000000110001110000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_B(60) <= "0000000000001110011100000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_B(61) <= "0000000000001110111000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_B(62) <= "0000000000001111110000000000000000000000000000000000000000000000";
SpaceShip_Frame_Fire_B(63) <= "0000000000001111100000000000000000000000000000000000000000000000";


-- Create integer versions of the row and column trackers
rowInt <= to_integer(unsigned(row));
colInt <= to_integer(unsigned(col));

-- VGA synchronisation block
uVGASync: VGASync
	port map(
		clk 	=> clk25,
		rst 	=> rst,
		hSync => hSync,
		vSync => vSync,
		row	=> row,
		col	=>	col,
		vidOn	=> vidOn
   );
  
-- Generate a 25Mhz clock from a 50MHz clock
ClkGen : process (clk50, rst)
begin
	if(rst = '0') then
		clk25 <= '0';
   elsif(clk50'event and clk50='1') then
    clk25 <= not(clk25);
	 clkCnt <= std_logic_vector(unsigned(clkCnt) + 1);
  end if;
end process;

clkTick <= clkCnt(23);
MovementTick <= clkCnt(17);
scoreTick <= clkCnt(18);

-- Track the pixel location and trace RGB values to the pixel
-- VGA Display 640 x 480: x is 0 -> 639, y is 0 -> 479
TraceXYPixels : process (clk25, rst, vidOn, rowInt, colInt, spaceShipX, score_Tracker1000, fireSignal, clkTick, alien1_X, alien1_Y, alien2_X, alien2_Y, alien3_X, alien3_Y, alien4_X, alien4_Y, alien5_X, alien5_Y)
variable x: integer :=0; -- Row pixel
variable y: integer :=0; -- Column pixel
variable c: integer :=0;
variable r: integer :=0;
variable offset128: integer := 127;
variable offset64: integer :=63;
variable offset32: integer :=31;
variable offset16: integer :=15;
variable offset8: integer :=7;
variable scoreOffset : integer := 120;
variable timeSwitch: boolean := false;
variable data: std_logic;

variable colour : std_logic_vector(2 downto 0);
begin
	-- Create variables from the input signals
	x := colInt;
	y := rowInt;
	if(clkTick'event and clkTick = '1') then
		if(timeSwitch = false) then
			timeSwitch := true;
		elsif(timeSwitch = true) then
			timeSwitch := false;
		else
			timeSwitch := false;
		end if;
	end if;
	-- If reset, set default RGB values (black)
	if(rst='0') then
		rgb <= "000";
	-- Otherwise, draw a pixel
	elsif(clk25'event and clk25 = '1') then
		if ((x >= scoreOffset) and (x <= scoreOffset+offset16) and (y >= 30) and (y <= 30+offset16)) then
		c := x - scoreOffset;
		r := y - 30;
		
		data := Score_S(r)(offset16-c);
		if(data = '1') then
			colour := "111";
		else
			colour := "000";
		end if;	
	elsif ((x >= scoreOffset+20) and (x <= scoreOffset+20+offset16) and (y >= 30) and (y <= 30+offset16)) then
		c := x - (scoreOffset+20);
		r := y - 30;
		
		data := Score_C(r)(offset16-c);
		if(data = '1') then
			colour := "111";
		else
			colour := "000";
		end if;	
	elsif ((x >= scoreOffset+40) and (x <= scoreOffset+40+offset16) and (y >= 30) and (y <= 30+offset16)) then
		c := x - (scoreOffset+40);
		r := y - 30;
		
		data := Score_O(r)(offset16-c);
		if(data = '1') then
			colour := "111";
		else
			colour := "000";
		end if;	
		elsif ((x >= scoreOffset+60) and (x <= scoreOffset+60+offset16) and (y >= 30) and (y <= 30+offset16)) then
			c := x - (scoreOffset+60);
			r := y - 30;
			
			data := Score_R(r)(offset16-c);
			if(data = '1') then
				colour := "111";
			else
				colour := "000";
			end if;
		elsif ((x >= scoreOffset+80) and (x <= scoreOffset+80+offset16) and (y >= 30) and (y <= 30+offset16)) then
			c := x - (scoreOffset+80);
			r := y - 30;
			
			data := Score_E(r)(offset16-c);
			if(data = '1') then
				colour := "111";
			else
				colour := "000";
			end if;
		elsif ((x >= scoreOffset+100) and (x <= scoreOffset+100+offset16) and (y >= 30) and (y <= 30+offset16)) then
			c := x - (scoreOffset+100);
			r := y - 30;
			
			data := Score_Semi(r)(offset16-c);
			if(data = '1') then
				colour := "111";
			else
				colour := "000";
			end if;
		elsif ((x >= scoreOffset+120) and (x <= scoreoffset+120+offset16) and (y >= 30) and (y <= 30+offset16)) then
			c := x - (scoreOffset+120);
			r := y - 30;
								
			data := Score_Tracker10000000000(r)(offset16-c);
			if(data = '1') then
				colour := "111";
			else
				colour := "000";
			end if;
		elsif ((x >= scoreOffset+140) and (x <= scoreoffset+140+offset16) and (y >= 30) and (y <= 30+offset16)) then
			c := x - (scoreOffset+140);
			r := y - 30;
								 
			data := Score_Tracker1000000000(r)(offset16-c);
			if(data = '1') then
				colour := "111";
			else
				colour := "000";
			end if;
		elsif ((x >= scoreOffset+160) and (x <= scoreoffset+160+offset16) and (y >= 30) and (y <= 30+offset16)) then
			c := x - (scoreOffset+160);
			r := y - 30;
								 
			data := Score_Tracker10000000(r)(offset16-c);
			if(data = '1') then
				colour := "111";
			else
				colour := "000";
			end if;
		elsif ((x >= scoreOffset+180) and (x <= scoreoffset+180+offset16) and (y >= 30) and (y <= 30+offset16)) then
			c := x - (scoreOffset+180);
			r := y - 30;
			
			data := Score_Tracker1000000(r)(offset16-c);
			if(data = '1') then
				colour := "111";
			else
				colour := "000";
			end if;
		elsif ((x >= scoreOffset+200) and (x <= scoreoffset+200+offset16) and (y >= 30) and (y <= 30+offset16)) then
			c := x - (scoreOffset+200);
			r := y - 30;
			
			data := Score_Tracker100000(r)(offset16-c);
			if(data = '1') then
				colour := "111";
			else
				colour := "000";
			end if;
		elsif ((x >= scoreOffset+220) and (x <= scoreoffset+220+offset16) and (y >= 30) and (y <= 30+offset16)) then
			c := x - (scoreOffset+220);
			r := y - 30;
			
			data := Score_Tracker10000(r)(offset16-c);
			if(data = '1') then
				colour := "111";
			else
				colour := "000";
			end if;
		elsif ((x >= scoreOffset+240) and (x <= scoreoffset+240+offset16) and (y >= 30) and (y <= 30+offset16)) then
			c := x - (scoreOffset+240);
			r := y - 30;
			
			data := Score_Tracker1000(r)(offset16-c);
			if(data = '1') then
				colour := "111";
			else
				colour := "000";
			end if;
		elsif ((x >= scoreOffset+260) and (x <= scoreOffset+260+offset16) and (y >= 30) and (y <= 30+offset16)) then
			c := x - (scoreOffset+260);
			r := y - 30;
			
			data := Score_Tracker100(r)(offset16-c);
			if(data = '1') then
				colour := "111";
			else
				colour := "000";
			end if;
		elsif ((x >= scoreOffset+280) and (x <= scoreOffset+280+offset16) and (y >= 30) and (y <= 30+offset16)) then
			c := x -  (scoreOffset+280);
			r := y - 30;
			
			data := Score_Tracker10(r)(offset16-c);
			if(data = '1') then
				colour := "111";
			else
				colour := "000";
			end if;
		elsif ((x >= scoreOffset+300) and (x <= scoreOffset+300+offset16) and (y >= 30) and (y <= 30+offset16)) then
			c := x - (scoreOffset+300);
			r := y - 30;
			
			data := Score_0(r)(offset16-c);
			if(data = '1') then
				colour := "111";
			else
				colour := "000";
			end if;
		elsif(gameOver = '0') then
			if((x >= 50) and (x <= 50+offset64) and (y >= spaceShipX-offset32) and (y <= spaceShipX+offset32) and (fireSignal = '1')) then
				c := x - 50;
				r := y - (spaceShipX-offset32);
				
				data := SpaceShip_Frame_Fire_R(r)(offset64-c);
				if(data = '1') then
					colour(2) := '1';
				else
					colour(2) := '0';
				end if;
				data := SpaceShip_Frame_Fire_G(r)(offset64-c);
				if(data = '1') then
					colour(1) := '1';
				else
					colour(1) := '0';
				end if;
				data := SpaceShip_Frame_Fire_B(r)(offset64-c);
				if(data = '1') then
					colour(0) := '1';
				else
					colour(0) := '0';
				end if;
				elsif((x >= 50) and (x <= 50+offset64) and (y >= spaceShipX-offset32) and (y <= spaceShipX+offset32) and (timeSwitch = false)) then
				c := x - 50;
				r := y - (spaceShipX-offset32);
				
				data := SpaceShip_Frame1_R(r)(offset64-c);
				if(data = '1') then
					colour(2) := '1';
				else
					colour(2) := '0';
				end if;
				data := SpaceShip_Frame1_G(r)(offset64-c);
				if(data = '1') then
					colour(1) := '1';
				else
					colour(1) := '0';
				end if;
				data := SpaceShip_Frame1_B(r)(offset64-c);
				if(data = '1') then
					colour(0) := '1';
				else
					colour(0) := '0';
				end if;
				elsif((x >= 50) and (x <= 50+offset64) and (y >= spaceShipX-offset32) and (y <= spaceShipX+offset32) and (timeSwitch = true)) then
				c := x - 50;
				r := y - (spaceShipX-offset32);
				
				data := SpaceShip_Frame2_R(r)(offset64-c);
				if(data = '1') then
					colour(2) := '1';
				else
					colour(2) := '0';
				end if;
				data := SpaceShip_Frame2_G(r)(offset64-c);
				if(data = '1') then
					colour(1) := '1';
				else
					colour(1) := '0';
				end if;
				data := SpaceShip_Frame2_B(r)(offset64-c);
				if(data = '1') then
					colour(0) := '1';
				else
					colour(0) := '0';
				end if;
				elsif((x >= bulletX) and (x<= bulletX+offset16) and (y >= bulletY-offset8) and (y <= bulletY+offset8) and timeSwitch = false) then
				if(fireSignal = '1') then
					c := x - BulletX;
					r := y - (BulletY + offset32 + offset8 + 4);
					
					data := Fire_Blast_1_R(r)(offset32-c);
					if(data = '1') then
						colour(2) := '1';
					else
						colour(2) := '0';
					end if;
					data := Fire_Blast_1_G(r)(offset32-c);
					if(data = '1') then
						colour(1) := '1';
					else
						colour(1) := '0';
					end if;
					data := Fire_Blast_1_B(r)(offset32-c);
					if(data = '1') then
						colour(0) := '1';
					else
						colour(0) := '0';
					end if;
				else
					colour := "000";
				end if;
				elsif((x >= bulletX) and (x<= bulletX+offset16) and (y >= bulletY-offset8) and (y <= bulletY+offset8) and timeSwitch = true) then
				if(fireSignal = '1') then
					c := x - BulletX;
					r := y - (BulletY + offset32 + offset8 + 4);
					
					data := Fire_Blast_2_R(r)(offset32-c);
					if(data = '1') then
						colour(2) := '1';
					else
						colour(2) := '0';
					end if;
					data := Fire_Blast_2_G(r)(offset32-c);
					if(data = '1') then
						colour(1) := '1';
					else
						colour(1) := '0';
					end if;
					data := Fire_Blast_2_B(r)(offset32-c);
					if(data = '1') then
						colour(0) := '1';
					else
						colour(0) := '0';
					end if;
				else
					colour := "000";
				end if;
				elsif((x >= Alien1_X) and (x<= Alien1_X+offset32) and (y >= Alien1_Y-offset16) and (y <= Alien1_Y+offset16) and timeSwitch = false and alien1_alive = '1') then
					c := x - Alien1_X;
					r := y - (Alien1_Y + offset16);
					
					data := Alien_1_R(r)(offset32-c);
					if(data = '1') then
						colour(2) := '1';
					else
						colour(2) := '0';
					end if;
					data := Alien_1_G(r)(offset32-c);
					if(data = '1') then
						colour(1) := '1';
					else
						colour(1) := '0';
					end if;
					data := Alien_1_B(r)(offset32-c);
					if(data = '1') then
						colour(0) := '1';
					else
						colour(0) := '0';
					end if;
			
				elsif((x >= Alien1_X) and (x<= Alien1_X+offset32) and (y >= Alien1_Y-offset16) and (y <= Alien1_Y+offset16) and timeSwitch = true and alien1_alive = '1') then
					c := x - Alien1_X;
					r := y - (Alien1_Y + offset16);
					
					data := Alien_2_R(r)(offset32-c);
					if(data = '1') then
						colour(2) := '1';
					else
						colour(2) := '0';
					end if;
					data := Alien_2_G(r)(offset32-c);
					if(data = '1') then
						colour(1) := '1';
					else
						colour(1) := '0';
					end if;
					data := Alien_2_B(r)(offset32-c);
					if(data = '1') then
						colour(0) := '1';
					else
						colour(0) := '0';
					end if;
				elsif((x >= Alien2_X) and (x<= Alien2_X+offset32) and (y >= Alien2_Y-offset16) and (y <= Alien2_Y+offset16) and timeSwitch = true and Alien2_alive = '1') then
					c := x - Alien2_X;
					r := y - (Alien2_Y + offset16);
					
					data := Alien_1_R(r)(offset32-c);
					if(data = '1') then
						colour(2) := '1';
					else
						colour(2) := '0';
					end if;
					data := Alien_1_G(r)(offset32-c);
					if(data = '1') then
						colour(1) := '1';
					else
						colour(1) := '0';
					end if;
					data := Alien_1_B(r)(offset32-c);
					if(data = '1') then
						colour(0) := '1';
					else
						colour(0) := '0';
					end if;
			
				elsif((x >= Alien2_X) and (x<= Alien2_X+offset32) and (y >= Alien2_Y-offset16) and (y <= Alien2_Y+offset16) and timeSwitch = false and Alien2_alive = '1') then
					c := x - Alien2_X;
					r := y - (Alien2_Y + offset16);
					
					data := Alien_2_R(r)(offset32-c);
					if(data = '1') then
						colour(2) := '1';
					else
						colour(2) := '0';
					end if;
					data := Alien_2_G(r)(offset32-c);
					if(data = '1') then
						colour(1) := '1';
					else
						colour(1) := '0';
					end if;
					data := Alien_2_B(r)(offset32-c);
					if(data = '1') then
						colour(0) := '1';
					else
						colour(0) := '0';
					end if;
				elsif((x >= Alien3_X) and (x<= Alien3_X+offset32) and (y >= Alien3_Y-offset16) and (y <= Alien3_Y+offset16) and timeSwitch = false and Alien3_alive = '1') then
					c := x - Alien3_X;
					r := y - (Alien3_Y + offset16);
					
					data := Alien_1_R(r)(offset32-c);
					if(data = '1') then
						colour(2) := '1';
					else
						colour(2) := '0';
					end if;
					data := Alien_1_G(r)(offset32-c);
					if(data = '1') then
						colour(1) := '1';
					else
						colour(1) := '0';
					end if;
					data := Alien_1_B(r)(offset32-c);
					if(data = '1') then
						colour(0) := '1';
					else
						colour(0) := '0';
					end if;
			
				elsif((x >= Alien3_X) and (x<= Alien3_X+offset32) and (y >= Alien3_Y-offset16) and (y <= Alien3_Y+offset16) and timeSwitch = true and Alien3_alive = '1') then
					c := x - Alien3_X;
					r := y - (Alien3_Y + offset16);
					
					data := Alien_2_R(r)(offset32-c);
					if(data = '1') then
						colour(2) := '1';
					else
						colour(2) := '0';
					end if;
					data := Alien_2_G(r)(offset32-c);
					if(data = '1') then
						colour(1) := '1';
					else
						colour(1) := '0';
					end if;
					data := Alien_2_B(r)(offset32-c);
					if(data = '1') then
						colour(0) := '1';
					else
						colour(0) := '0';
					end if;
				elsif((x >= Alien4_X) and (x<= Alien4_X+offset32) and (y >= Alien4_Y-offset16) and (y <= Alien4_Y+offset16) and timeSwitch = true and Alien4_alive = '1') then
					c := x - Alien4_X;
					r := y - (Alien4_Y + offset16);
					
					data := Alien_1_R(r)(offset32-c);
					if(data = '1') then
						colour(2) := '1';
					else
						colour(2) := '0';
					end if;
					data := Alien_1_G(r)(offset32-c);
					if(data = '1') then
						colour(1) := '1';
					else
						colour(1) := '0';
					end if;
					data := Alien_1_B(r)(offset32-c);
					if(data = '1') then
						colour(0) := '1';
					else
						colour(0) := '0';
					end if;
			
				elsif((x >= Alien4_X) and (x<= Alien4_X+offset32) and (y >= Alien4_Y-offset16) and (y <= Alien4_Y+offset16) and timeSwitch = false and Alien4_alive = '1') then
					c := x - Alien4_X;
					r := y - (Alien4_Y + offset16);
					
					data := Alien_2_R(r)(offset32-c);
					if(data = '1') then
						colour(2) := '1';
					else
						colour(2) := '0';
					end if;
					data := Alien_2_G(r)(offset32-c);
					if(data = '1') then
						colour(1) := '1';
					else
						colour(1) := '0';
					end if;
					data := Alien_2_B(r)(offset32-c);
					if(data = '1') then
						colour(0) := '1';
					else
						colour(0) := '0';
					end if;
				elsif((x >= Alien5_X) and (x<= Alien5_X+offset32) and (y >= Alien5_Y-offset16) and (y <= Alien5_Y+offset16) and timeSwitch = false and Alien5_alive = '1') then
					c := x - Alien5_X;
					r := y - (Alien5_Y + offset16);
					
					data := Alien_1_R(r)(offset32-c);
					if(data = '1') then
						colour(2) := '1';
					else
						colour(2) := '0';
					end if;
					data := Alien_1_G(r)(offset32-c);
					if(data = '1') then
						colour(1) := '1';
					else
						colour(1) := '0';
					end if;
					data := Alien_1_B(r)(offset32-c);
					if(data = '1') then
						colour(0) := '1';
					else
						colour(0) := '0';
					end if;
			
				elsif((x >= Alien5_X) and (x<= Alien5_X+offset32) and (y >= Alien5_Y-offset16) and (y <= Alien5_Y+offset16) and timeSwitch = true and Alien5_alive = '1') then
					c := x - Alien5_X;
					r := y - (Alien5_Y + offset16);
					
					data := Alien_2_R(r)(offset32-c);
					if(data = '1') then
						colour(2) := '1';
					else
						colour(2) := '0';
					end if;
					data := Alien_2_G(r)(offset32-c);
					if(data = '1') then
						colour(1) := '1';
					else
						colour(1) := '0';
					end if;
					data := Alien_2_B(r)(offset32-c);
					if(data = '1') then
						colour(0) := '1';
					else
						colour(0) := '0';
					end if;
				else
				colour := "000";
				end if;
		elsif(gameOver = '1') then
			if ((x >= 250) and (x <= 250+offset16) and (y >= 220) and (y <= 220+offset16)) then
			c := x - 250;
			r := y - 220;
			
			data := GameOver_G_W(r)(offset16-c);
			if(data = '1') then
				colour := "111";
			else
				colour := "000";
			end if;
			elsif ((x >= 270) and (x <= 270+offset16) and (y >= 220) and (y <= 220+offset16)) then
			c := x - 270;
			r := y - 220;
			
			data := GameOver_A_W(r)(offset16-c);
			if(data = '1') then
				colour := "111";
			else
				colour := "000";
			end if;
			elsif ((x >= 290) and (x <= 290+offset16) and (y >= 220) and (y <= 220+offset16)) then
			c := x - 290;
			r := y - 220;
			
			data := GameOver_M_W(r)(offset16-c);
			if(data = '1') then
				colour := "111";
			else
				colour := "000";
			end if;
			elsif ((x >= 310) and (x <= 310+offset16) and (y >= 220) and (y <= 220+offset16)) then
			c := x - 310;
			r := y - 220;
			
			data := Score_E(r)(offset16-c);
			if(data = '1') then
				colour := "111";
			else
				colour := "000";
			end if;
			elsif ((x >= 340) and (x <= 340+offset16) and (y >= 220) and (y <= 220+offset16)) then
			c := x - 340;
			r := y - 220;
			
			data := Score_O(r)(offset16-c);
			if(data = '1') then
				colour := "111";
			else
				colour := "000";
			end if;
			elsif ((x >= 360) and (x <= 360+offset16) and (y >= 220) and (y <= 220+offset16)) then
			c := x - 360;
			r := y - 220;
			
			data := GameOver_V_W(r)(offset16-c);
			if(data = '1') then
				colour := "111";
			else
				colour := "000";
			end if;
		elsif ((x >= 380) and (x <= 380+offset16) and (y >= 220) and (y <= 220+offset16)) then
			c := x - 380;
			r := y - 220;
			
			data := Score_E(r)(offset16-c);
			if(data = '1') then
				colour := "111";
			else
				colour := "000";
			end if;
		elsif ((x >= 400) and (x <= 400+offset16) and (y >= 220) and (y <= 220+offset16)) then
			c := x - 400;
			r := y - 220;
			
			data := Score_R(r)(offset16-c);
			if(data = '1') then
				colour := "111";
			else
				colour := "000";
			end if;
		else 
			colour := "000";
		end if;
	
		end if;
		rgb <= colour;
	end if;
end process;

StarShipMovement:process(movementTick, rst, downButton, upButton, startDebounce, clk50, rotary_event, rotary_left)
variable y: integer :=320; 
begin
	if(rst = '0') then
		y := 320;
	elsif(clk50'event and	clk50 = '1') then
		if(rotary_event = '1' and rotary_left = '0') then
				y := y + 5;
				if(y >= 440) then 
					y := 440;
				end if;
		elsif(rotary_event = '1' and rotary_left = '1') then
				y := y - 5;
				if(y <= 100) then 
					y := 100;
				end if;
		end if;

		

		spaceShipX <= y;
	end if;
end process;



gameOverSwitch:Process(movementTick, rst, spaceshipX, alien1_X, alien1_Y, alien2_X, alien2_Y, alien3_X, alien3_Y, alien4_X, alien4_Y, alien5_X, alien5_Y)
begin
	if(rst = '0') then
		gameOver <= '0';
	elsif(movementTick'event and movementTick = '1') then
			if(alien1_Y >= (spaceshipX-32) and alien1_Y <= (spaceshipX+32) and alien1_X <= 100) then
					gameOver <= '1';
			elsif(alien2_Y >= (spaceshipX-32) and alien2_Y <= (spaceshipX+32) and alien2_X <= 100) then
					gameOver <= '1';
			elsif(alien3_Y >= (spaceshipX-32) and alien3_Y <= (spaceshipX+32) and alien3_X <= 100) then
					gameOver <= '1';
			elsif (alien4_Y >= (spaceshipX-32) and alien4_Y <= (spaceshipX+32) and alien4_X <= 100) then
					gameOver <= '1';
			elsif(alien5_Y >= (spaceshipX-32) and alien5_Y <= (spaceshipX+32) and alien5_X <= 100) then
					gameOver <= '1';
			end if;
	end if;
end process;

alien1Alive:process(movementTick, rst)
variable alive : std_logic := '0';
begin
	if(rst = '0') then
		alive := '0';
	elsif(movementTick'event and	movementTick = '1') then
		if(BulletX >= alien1_X and BulletX <= alien1_X+32 and BulletY >= alien1_Y-16 and BulletY <= alien1_Y+16) then
			alive := '0';
		elsif(alien1_X >= 540) then
			alive := '1';
		end if; 
		alien1_alive <= alive;
	end if;
end process;

alien1Movement:process(clkTick, rst, SpaceshipX, alien1_alive)
variable y: integer :=116; 
variable x: integer :=560;
begin
	if(rst = '0') then
		y := 116;
		x := 560;
	elsif(clkTick'event and	clkTick = '1') then
		if(x >= 50) then
			x := x - 26;
		else
			if( y < SpaceshipX ) then
					y := y + 5;
			elsif( y > SpaceshipX ) then
					y := y - 5;
			end if;
		end if;
		if(alien1_alive = '0') then
			x := 560;
			y := 116;
		end if;
		alien1_Y <= y;
		alien1_X <= x;
	end if;
end process;

alien2Alive:process(movementTick, rst, SpaceshipX, alien2_alive)
variable alive : std_logic := '0';
begin
	if(rst = '0') then
		alive := '0';
	elsif(movementTick'event and	movementTick = '1') then
		if(BulletX >= alien2_X and BulletX <= alien2_X+32 and BulletY >= alien2_Y-16 and BulletY <= alien2_Y+16) then
			alive := '0';
		elsif(alien2_X >= 540) then
			alive := '1';
		end if; 
		alien2_alive <= alive;
	end if;
end process;

alien2Movement:process(clkTick, rst, SpaceshipX, alien2_alive)
variable y: integer :=266; 
variable x: integer :=560;
begin
	if(rst = '0') then
		y := 266;
	x := 560;
	elsif(clkTick'event and	clkTick = '1') then
		if(x >= 50) then
			x := x - 24;
		else
			if( y < SpaceshipX ) then
					y := y + 5;
			elsif( y > SpaceshipX ) then
					y := y - 5;
			end if;
		end if;
		if(alien2_alive = '0') then
			x := 560;
			y := 266;
		end if;
		alien2_Y <= y;
		alien2_X <= x;
	end if;
end process;

alien3Alive:process(movementTick, rst, SpaceshipX, alien3_alive)
variable alive : std_logic := '0';
begin
	if(rst = '0') then
		alive := '0';
	elsif(movementTick'event and	movementTick = '1') then
		if(BulletX >= alien3_X and BulletX <= alien3_X+32 and BulletY >= alien3_Y-16 and BulletY <= alien3_Y+16) then
			alive := '0';
		elsif(alien3_X >= 540) then
			alive := '1';
		end if; 
		alien3_alive <= alive;
	end if;
end process;

alien3Movement:process(clkTick, rst, SpaceshipX, alien3_alive)
variable y: integer :=416; 
variable x: integer :=560;
begin
	if(rst = '0') then
		y := 416;
	x := 560;
	elsif(clkTick'event and	clkTick = '1') then
		if(x >= 50) then
			x := x - 20;
		else
			if( y < SpaceshipX ) then
					y := y + 5;
			elsif( y > SpaceshipX ) then
					y := y - 5;
			end if;
		end if;
		if(alien3_alive = '0') then
			x := 560;
			y := 416;
		end if;
		alien3_Y <= y;
		alien3_X <= x;
	end if;
end process;

alien4Alive:process(movementTick, rst)
variable alive : std_logic := '0';
begin
	if(rst = '0') then
		alive := '0';
	elsif(movementTick'event and	movementTick = '1') then
		if(BulletX >= alien4_X and BulletX <= alien4_X+32 and BulletY >= alien4_Y-16 and BulletY <= alien4_Y+16) then
			alive := '0';
		elsif(alien4_X >= 540) then
			alive := '1';
		end if; 
		alien4_alive <= alive;
	end if;
end process;

alien4Movement:process(clkTick, rst)
variable y: integer :=316; 
variable x: integer :=560;
begin
	if(rst = '0') then
		y := 316;
		x := 560;
	elsif(clkTick'event and	clkTick = '1') then
		if(x >= 50) then
			x := x - 21;
		else
			if( y < SpaceshipX ) then
					y := y + 5;
			elsif( y > SpaceshipX ) then
					y := y - 5;
			end if;
		end if;
		if(alien4_alive = '0') then
			x := 560;
			y := 316;
		end if;
		alien4_Y <= y;
		alien4_X <= x;
	end if;
end process;

alien5Alive:process(movementTick, rst)
variable alive : std_logic := '0';
begin
	if(rst = '0') then
		alive := '0';
	elsif(movementTick'event and	movementTick = '1') then
		if(BulletX >= alien5_X and BulletX <= alien5_X+32 and BulletY >= alien5_Y-16 and BulletY <= alien5_Y+16) then
			alive := '0';
		elsif(alien5_X >= 540) then
			alive := '1';
		end if; 
		alien5_alive <= alive;
	end if;
end process;

alien5Movement:process(clkTick, rst)
variable y: integer :=216; 
variable x: integer :=560;
begin
	if(rst = '0') then
		y := 216;
	x := 560;
	elsif(clkTick'event and	clkTick = '1') then
		if(x >= 50) then
			x := x - 25;
		else
			if( y < SpaceshipX ) then
					y := y + 5;
			elsif( y > SpaceshipX ) then
					y := y - 5;
			end if;
		end if;
		if(alien5_alive = '0') then
			x := 560;
			y := 216;
		end if;
		alien5_Y <= y;
		alien5_X <= x;
	end if;
end process;

SpaceShipShoot:process(movementTick, rst, fireButton)
variable fireTemp : std_logic := '0';
begin
	if(rst = '0') then
		fireTemp := '0';
	elsif(movementTick'event and movementTick = '1') then
		if(fireButton = '1') then
			fireTemp := '1';
		elsif(fireButton = '0' and BulletX >= 620) then 
			fireTemp := '0';
		end if;
	end if;
	fireSignal <= fireTemp;
end process;

fireAnimation:process(rst, movementTick, spaceShipX, fireSignal)
	variable x : integer range 114 to 630;
	variable y : integer := 0;
	variable fired : boolean := false;
begin
	if(rst = '0') then 
		bulletX <= 114;
		bulletY <= spaceShipX;
		x := 114;
		y := spaceShipX;
	elsif(movementTick'event and movementTick = '1') then
		if(fireSignal = '1' and startDebounce = true and fired = false) then 
			fired := true;
			y := SpaceshipX;
		end if;
		if(fired = true) then
			BulletY <= y;
				x := x+5;
				if(x >= 630) then
					fired := false;
					x := 114; 
				end if; 
		end if;
		BulletX <= x;
		BulletY <= y;
	end if;
end process;




CalcScore:process(rst, scoreTick, score10, score100, score1000, alien1_alive, alien2_alive, alien3_alive, alien4_alive, alien5_alive)

	variable scoreTemp : integer := 0;
begin
	if(rst = '0') then 
			score1000000000 <= 0;
			score100000000 <= 0;
			score10000000 <= 0; 
			score1000000 <= 0;
			score100000 <= 0; 
			score10000 <= 0;
			score1000 <= 0; 
			score100 <= 0;
			score10 <= 0; 
	else
		if(scoreTick'event and scoreTick = '1') then 
			if(alien1_alive = '0' or alien2_alive = '0' or alien3_alive = '0' or alien4_alive = '0' or alien5_alive = '0') then
				score10 <= score10+1;
				if(score10 = 10) then
					score10 <= 0; 
					score100 <= score100 + 1;
					if(score100 = 10) then
						score1000 <= score1000 + 1;
						score100 <= 0;
						if(score1000 = 10) then
							score1000 <= 0;
							score10000 <= score10000 + 1;
							if(score10000 = 10) then
								score10000 <= 0; 
								score100000 <= score100000 + 1;
								if(score100000 = 10) then
									score100000 <= 0;
									score1000000 <= score1000000 + 1;
									if(score1000000 = 10) then
										score1000000 <= 0;
										score10000000 <= score10000000 + 1;
										if(score10000000 = 10) then
											score10000000 <= 0;
											score100000000 <= score100000000 + 1;
											if(score100000000 = 10) then
												score100000000 <= 0;
												score1000000000 <= score1000000000 + 1;
												if(score1000000000 = 10) then
													score1000000000 <= 0;
													score10000000000 <= score10000000000 + 1;
												end if;
											end if;
										end if;
									end if;
								end if;
							end if;
						end if;
					end if;
				end if;
			end if;
		end if;
	end if;
end process;

DisplayScore: process(clkTick, rst, score10, score100, score1000)
begin
	if(rst = '0') then
		for I in 0 to 15 loop
			Score_Tracker10000000000(I) <= "0000000000000000";
			Score_Tracker1000000000(I) <= "0000000000000000";
			Score_Tracker100000000(I) <= "0000000000000000";
			Score_Tracker10000000(I) <= "0000000000000000";
			Score_Tracker1000000(I) <= "0000000000000000";
			Score_Tracker100000(I) <= "0000000000000000";
			Score_Tracker10000(I) <= "0000000000000000";
			Score_Tracker1000(I) <= "0000000000000000";
			Score_Tracker100(I) <= "0000000000000000";
			Score_Tracker10(I) <= "0000000000000000";
		end loop;
	elsif(clkTick'event and clkTick = '1') then 
	if(score10000000000 = 0) then
			Score_Tracker10000000000 <= Score_0;
		elsif(score10000000000 = 1) then
			Score_Tracker10000000000 <= Score_1;
		elsif(score10000000000 = 2) then
			Score_Tracker10000000000 <= Score_2;
		elsif(score10000000000 = 3) then
			Score_Tracker10000000000 <= Score_3;
		elsif(score10000000000 = 4) then
			Score_Tracker10000000000 <= Score_4;
		elsif(score10000000000 = 5) then
			Score_Tracker10000000000 <= Score_5;
		elsif(score10000000000 = 6) then
			Score_Tracker10000000000 <= Score_6;
		elsif(score10000000000 = 7) then
			Score_Tracker10000000000 <= Score_7;
		elsif(score10000000000 = 8) then
			Score_Tracker10000000000 <= Score_8;
		elsif(score10000000000 = 9) then
			Score_Tracker10000000000 <= Score_9;
		end if;
	if(score1000000000 = 0) then
			Score_Tracker1000000000 <= Score_0;
		elsif(score1000000000 = 1) then
			Score_Tracker1000000000 <= Score_1;
		elsif(score1000000000 = 2) then
			Score_Tracker1000000000 <= Score_2;
		elsif(score1000000000 = 3) then
			Score_Tracker1000000000 <= Score_3;
		elsif(score1000000000 = 4) then
			Score_Tracker1000000000 <= Score_4;
		elsif(score1000000000 = 5) then
			Score_Tracker1000000000 <= Score_5;
		elsif(score1000000000 = 6) then
			Score_Tracker1000000000 <= Score_6;
		elsif(score1000000000 = 7) then
			Score_Tracker1000000000 <= Score_7;
		elsif(score1000000000 = 8) then
			Score_Tracker1000000000 <= Score_8;
		elsif(score1000000000 = 9) then
			Score_Tracker1000000000 <= Score_9;
		end if;
	if(score100000000 = 0) then
			Score_Tracker100000000 <= Score_0;
		elsif(score100000000 = 1) then
			Score_Tracker100000000 <= Score_1;
		elsif(score100000000 = 2) then
			Score_Tracker100000000 <= Score_2;
		elsif(score100000000 = 3) then
			Score_Tracker100000000 <= Score_3;
		elsif(score100000000 = 4) then
			Score_Tracker100000000 <= Score_4;
		elsif(score100000000 = 5) then
			Score_Tracker100000000 <= Score_5;
		elsif(score100000000 = 6) then
			Score_Tracker100000000 <= Score_6;
		elsif(score100000000 = 7) then
			Score_Tracker100000000 <= Score_7;
		elsif(score100000000 = 8) then
			Score_Tracker100000000 <= Score_8;
		elsif(score100000000 = 9) then
			Score_Tracker100000000 <= Score_9;
		end if;
	if(score10000000 = 0) then
			Score_Tracker10000000 <= Score_0;
		elsif(score10000000 = 1) then
			Score_Tracker10000000 <= Score_1;
		elsif(score10000000 = 2) then
			Score_Tracker10000000 <= Score_2;
		elsif(score10000000 = 3) then
			Score_Tracker10000000 <= Score_3;
		elsif(score10000000 = 4) then
			Score_Tracker10000000 <= Score_4;
		elsif(score10000000 = 5) then
			Score_Tracker10000000 <= Score_5;
		elsif(score10000000 = 6) then
			Score_Tracker10000000 <= Score_6;
		elsif(score10000000 = 7) then
			Score_Tracker10000000 <= Score_7;
		elsif(score10000000 = 8) then
			Score_Tracker10000000 <= Score_8;
		elsif(score10000000 = 9) then
			Score_Tracker10000000 <= Score_9;
		end if;
	if(score1000000 = 0) then
			Score_Tracker1000000 <= Score_0;
		elsif(score1000000 = 1) then
			Score_Tracker1000000 <= Score_1;
		elsif(score1000000 = 2) then
			Score_Tracker1000000 <= Score_2;
		elsif(score1000000 = 3) then
			Score_Tracker1000000 <= Score_3;
		elsif(score1000000 = 4) then
			Score_Tracker1000000 <= Score_4;
		elsif(score1000000 = 5) then
			Score_Tracker1000000 <= Score_5;
		elsif(score1000000 = 6) then
			Score_Tracker1000000 <= Score_6;
		elsif(score1000000 = 7) then
			Score_Tracker1000000 <= Score_7;
		elsif(score1000000 = 8) then
			Score_Tracker1000000 <= Score_8;
		elsif(score1000000 = 9) then
			Score_Tracker1000000 <= Score_9;
		end if;
	
		if(score100000 = 0) then
			Score_Tracker100000 <= Score_0;
		elsif(score100000 = 1) then
			Score_Tracker100000 <= Score_1;
		elsif(score100000 = 2) then
			Score_Tracker100000 <= Score_2;
		elsif(score100000 = 3) then
			Score_Tracker100000 <= Score_3;
		elsif(score100000 = 4) then
			Score_Tracker100000 <= Score_4;
		elsif(score100000 = 5) then
			Score_Tracker100000 <= Score_5;
		elsif(score100000 = 6) then
			Score_Tracker100000 <= Score_6;
		elsif(score100000 = 7) then
			Score_Tracker100000 <= Score_7;
		elsif(score100000 = 8) then
			Score_Tracker100000 <= Score_8;
		elsif(score100000 = 9) then
			Score_Tracker100000 <= Score_9;
		end if;
		
		if(score10000 = 0) then
			Score_Tracker10000 <= Score_0;
		elsif(score10000 = 1) then
			Score_Tracker10000 <= Score_1;
		elsif(score10000 = 2) then
			Score_Tracker10000 <= Score_2;
		elsif(score10000 = 3) then
			Score_Tracker10000 <= Score_3;
		elsif(score10000 = 4) then
			Score_Tracker10000 <= Score_4;
		elsif(score10000 = 5) then
			Score_Tracker10000 <= Score_5;
		elsif(score10000 = 6) then
			Score_Tracker10000 <= Score_6;
		elsif(score10000 = 7) then
			Score_Tracker10000 <= Score_7;
		elsif(score10000 = 8) then
			Score_Tracker10000 <= Score_8;
		elsif(score10000 = 9) then
			Score_Tracker10000 <= Score_9;
		end if;
		if(score1000 = 0) then
			Score_Tracker1000 <= Score_0;
		elsif(score1000 = 1) then
			Score_Tracker1000 <= Score_1;
		elsif(score1000 = 2) then
			Score_Tracker1000 <= Score_2;
		elsif(score1000 = 3) then
			Score_Tracker1000 <= Score_3;
		elsif(score1000 = 4) then
			Score_Tracker1000 <= Score_4;
		elsif(score1000 = 5) then
			Score_Tracker1000 <= Score_5;
		elsif(score1000 = 6) then
			Score_Tracker1000 <= Score_6;
		elsif(score1000 = 7) then
			Score_Tracker1000 <= Score_7;
		elsif(score1000 = 8) then
			Score_Tracker1000 <= Score_8;
		elsif(score1000 = 9) then
			Score_Tracker1000 <= Score_9;
		end if;
		if(score100 = 0) then
			Score_Tracker100 <= Score_0;
		elsif(score100 = 1) then
			Score_Tracker100 <= Score_1;
		elsif(score100 = 2) then
			Score_Tracker100 <= Score_2;
		elsif(score100 = 3) then
			Score_Tracker100 <= Score_3;
		elsif(score100 = 4) then
			Score_Tracker100 <= Score_4;
		elsif(score100 = 5) then
			Score_Tracker100 <= Score_5;
		elsif(score100 = 6) then
			Score_Tracker100 <= Score_6;
		elsif(score100 = 7) then
			Score_Tracker100 <= Score_7;
		elsif(score100 = 8) then
			Score_Tracker100 <= Score_8;
		elsif(score100 = 9) then
			Score_Tracker100 <= Score_9;
		end if;
		if(score10 = 0) then
			Score_Tracker10 <= Score_0;
		elsif(score10 = 1) then
			Score_Tracker10 <= Score_1;
		elsif(score10 = 2) then
			Score_Tracker10 <= Score_2;
		elsif(score10 = 3) then
			Score_Tracker10 <= Score_3;
		elsif(score10 = 4) then
			Score_Tracker10 <= Score_4;
		elsif(score10 = 5) then
			Score_Tracker10 <= Score_5;
		elsif(score10 = 6) then
			Score_Tracker10 <= Score_6;
		elsif(score10 = 7) then
			Score_Tracker10 <= Score_7;
		elsif(score10 = 8) then
			Score_Tracker10 <= Score_8;
		elsif(score10 = 9) then
			Score_Tracker10 <= Score_9;
		end if;
	end if;
end process;
		
		
Debounce:process(rst, movementTick, startDebounce, debounceCounter, downButton, upButton, fireButton)
  begin
	if(rst = '0') then
		debounceCounter <= "1000";
	elsif (movementTick'event and movementTick = '1') then 
		if(startDebounce = false) then
			if ((downButton = '1') or (upButton = '1') or (fireButton = '1')) then
			  startDebounce <= true;
			end if;
		end if;

		if(startDebounce = true) then
			debounceCounter <= std_logic_vector(unsigned(debounceCounter) - 1);  
			if(debounceCounter = "1000") then
				debounceCounter <= "1000";
				startDebounce <= false;
			end if;
      end if;   
	end if;
end process;

rotary_filter: process(clk50, rotary_in, rotary_b_in, rotary_a_in)
begin
	if clk50'event and clk50='1' then
		rotary_in <= rotary_b_in & rotary_a_in;
		case rotary_in is
			when "00" =>
				rotary_q1 <= '0';
				rotary_q2 <= rotary_q2;
			when "01" => 
				rotary_q1 <= rotary_q1;
				rotary_q2 <= '0';
			when "10" => 
				rotary_q1 <= rotary_q1;
				rotary_q2 <= '1';
			when "11" => 
				rotary_q1 <= '1';
				rotary_q2 <= rotary_q2;
			when others => rotary_q1 <= rotary_q1;
				rotary_q2 <= rotary_q2;
		end case;
	end if;
end process rotary_filter;

direction: process(clk50)
begin
	if clk50'event and clk50='1' then
		delay_rotary_q1 <= rotary_q1;
		if rotary_q1='1' and delay_rotary_q1='0' then
			rotary_event <= '1';
			rotary_left <= rotary_q2;
		else
			rotary_event <= '0';
			rotary_left <= rotary_left;
		end if;
	end if;
end process direction;


-- Drive outputs
r <= rgb(2) and vidOn;
g <= rgb(1) and vidOn;
b <= rgb(0) and vidOn;

end RTL;


